#******
# TECH LIB NAME: smic18
# TECH FILE NAME: techfile.cds
#
# RC values have been extracted from SMIC's Interconnect Capacitance
# Table, Rev 2.0, Date 02-08-2003 and Document TD-L018-BL-2001 Rev 2R
#
# Resistance and Capacitance Values
# ---------------------------------
# The LEF technology files included in this directory contain
# resistance and capacitance (RC) values for the purpose of timing
# driven place & route.  Please note that the RC values contained in
# this tech file were created using the worst case interconnect models
# from the foundry and assume a full metal route at every grid location
# on every metal layer, so the values are intentionally very
# conservative. It is assumed that this technology file will be used
# only as a starting point for creating initial timing driven place &
# route runs during the development of your own more accurate RC
# values, tailored to your specific place & route environment. AS A
# RESULT, TIMING NUMBERS DERIVED FROM THESE RC VALUES MAY BE
# SIGNIFICANTLY SLOWER THAN REALITY.
#
# The RC values used in the LEF technology file are to be used only
# for timing driven place & route. Due to accuracy limitations,
# please do not attempt to use this file for chip-level RC extraction
# in conjunction with your sign-off timing simulations. For chip-level
# extraction, please use a dedicated extraction tool such as HyperExtract,
# starRC or Simplex, etc.
#
# $Id: smic18_6lm.lef,v 1.4 2003-03-10 18:30:04-08 wching Exp $
#
#******                                                               

VERSION 5.2 ;

NAMESCASESENSITIVE ON ;

UNITS
    DATABASE MICRONS 2000  ;
END UNITS

LAYER POLY1
    TYPE MASTERSLICE ;
END POLY1

LAYER METAL1
    TYPE ROUTING ;
    WIDTH 0.230 ;
    SPACING 0.230 ;
    SPACING 0.6 RANGE 10.0 100000.0 ;
    PITCH 0.560 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ      7.8000e-02 ;
    CAPACITANCE CPERSQDIST 1.1152e-04 ;
    EDGECAPACITANCE        9.0179e-05 ;
END METAL1

LAYER VIA12
    TYPE CUT ;
END VIA12

LAYER METAL2
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.6 RANGE 10.0 100000.0 ;
    PITCH 0.660 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ      7.8000e-02 ;
    CAPACITANCE CPERSQDIST 6.5875e-05 ;
    EDGECAPACITANCE        8.7917e-05 ;
END METAL2

LAYER VIA23
    TYPE CUT ;
END VIA23

LAYER METAL3
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.6 RANGE 10.0 100000.0 ;
    PITCH 0.560 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ      7.8000e-02 ;
    CAPACITANCE CPERSQDIST 5.9699e-05 ;
    EDGECAPACITANCE        1.0642e-04 ;
END METAL3

LAYER VIA34
    TYPE CUT ;
END VIA34

LAYER METAL4
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.6 RANGE 10.0 100000.0 ;
    PITCH 0.660 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ      7.8000e-02 ;
    CAPACITANCE CPERSQDIST 5.5911e-05 ;
    EDGECAPACITANCE        8.7491e-05 ;
END METAL4

LAYER VIA45
    TYPE CUT ;
END VIA45

LAYER METAL5
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.6 RANGE 10.0 100000.0 ;
    PITCH 1.120 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ      7.8000e-02 ;
    CAPACITANCE CPERSQDIST 4.3064e-05 ;
    EDGECAPACITANCE        5.6324e-05 ;
END METAL5

LAYER VIA56
    TYPE CUT ;
END VIA56

LAYER METAL6
    TYPE ROUTING ;
    WIDTH 0.440 ;
    SPACING 0.460 ;
    SPACING 0.6 RANGE 10.0 100000.0 ;
    PITCH 1.320 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ      3.6000e-02 ;
    CAPACITANCE CPERSQDIST 2.1886e-05 ;
    EDGECAPACITANCE        7.8084e-05 ;
END METAL6

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA via1 DEFAULT
    RESISTANCE 5.0000e+00 ;
    LAYER METAL1 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL2 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via1

VIA via2 DEFAULT
    RESISTANCE 5.0000e+00 ;
    LAYER METAL2 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via2

VIA via2ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 5.0000e+00 ;
    LAYER METAL2 ;
        RECT -0.140 -0.370 0.140 0.370 ;
    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via2ts

VIA via3 DEFAULT
    RESISTANCE 5.0000e+00 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL4 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via3

VIA via3ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 5.0000e+00 ;
    LAYER METAL3 ;
        RECT -0.370 -0.140 0.370 0.140 ;
    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL4 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via3ts

VIA via4 DEFAULT
    RESISTANCE 5.0000e+00 ;
    LAYER METAL4 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL5 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via4

VIA via4ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 5.0000e+00 ;
    LAYER METAL4 ;
        RECT -0.140 -0.370 0.140 0.370 ;
    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL5 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END via4ts

VIA via5 DEFAULT
    RESISTANCE 3.0000e+00 ;
    LAYER METAL5 ;
        RECT -0.240 -0.190 0.240 0.190 ;
    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METAL6 ;
        RECT -0.270 -0.270 0.270 0.270 ;
END via5

VIA via5ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 3.0000e+00 ;
    LAYER METAL5 ;
        RECT -0.270 -0.190 0.270 0.190 ;
    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METAL6 ;
        RECT -0.270 -0.270 0.270 0.270 ;
END via5ts

VIARULE via1Array GENERATE
    LAYER METAL1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER METAL2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END via1Array

VIARULE via2Array GENERATE
    LAYER METAL2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END via2Array

VIARULE via3Array GENERATE
    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER METAL4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END via3Array

VIARULE via4Array GENERATE
    LAYER METAL4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END via4Array

VIARULE via5Array GENERATE
    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER METAL6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
        SPACING 0.710 BY 0.710 ;
END via5Array

VIARULE TURNM1 GENERATE
    LAYER METAL1 ;
        DIRECTION vertical ;

    LAYER METAL1 ;
        DIRECTION horizontal ;
END TURNM1

VIARULE TURNM2 GENERATE
    LAYER METAL2 ;
        DIRECTION vertical ;

    LAYER METAL2 ;
        DIRECTION horizontal ;
END TURNM2

VIARULE TURNM3 GENERATE
    LAYER METAL3 ;
        DIRECTION vertical ;

    LAYER METAL3 ;
        DIRECTION horizontal ;
END TURNM3

VIARULE TURNM4 GENERATE
    LAYER METAL4 ;
        DIRECTION vertical ;

    LAYER METAL4 ;
        DIRECTION horizontal ;
END TURNM4

VIARULE TURNM5 GENERATE
    LAYER METAL5 ;
        DIRECTION vertical ;

    LAYER METAL5 ;
        DIRECTION horizontal ;
END TURNM5

VIARULE TURNM6 GENERATE
    LAYER METAL6 ;
        DIRECTION vertical ;

    LAYER METAL6 ;
        DIRECTION horizontal ;
END TURNM6

SPACING
    SAMENET METAL1 METAL1 0.230  ;
    SAMENET METAL2 METAL2 0.280 STACK ;
    SAMENET METAL3 METAL3 0.280 STACK ;
    SAMENET METAL4 METAL4 0.280 STACK ;
    SAMENET METAL5 METAL5 0.280 STACK ;
    SAMENET METAL6 METAL6 0.460  ;
    SAMENET VIA12 VIA12 0.260  ;
    SAMENET VIA23 VIA23 0.260  ;
    SAMENET VIA34 VIA34 0.260  ;
    SAMENET VIA45 VIA45 0.260  ;
    SAMENET VIA56 VIA56 0.350  ;
    SAMENET VIA12 VIA23 0.0 STACK ;
    SAMENET VIA23 VIA34 0.0 STACK ;
    SAMENET VIA34 VIA45 0.0 STACK ;
    SAMENET VIA45 VIA56 0.0 STACK ;
END SPACING

SITE smic18site
    SYMMETRY y  ;
    CLASS core  ;
    SIZE 0.660 BY 5.040 ;
END smic18site

MACRO FILL8
    CLASS CORE ;
    FOREIGN FILL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 5.280 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 5.280 5.440 ;
        END
    END VDD
END FILL8

MACRO FILL64
    CLASS CORE ;
    FOREIGN FILL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 42.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 42.240 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 42.240 5.440 ;
        END
    END VDD
END FILL64

MACRO FILL4
    CLASS CORE ;
    FOREIGN FILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 2.640 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 2.640 5.440 ;
        END
    END VDD
END FILL4

MACRO FILL32
    CLASS CORE ;
    FOREIGN FILL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 21.120 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 21.120 5.440 ;
        END
    END VDD
END FILL32

MACRO FILL2
    CLASS CORE ;
    FOREIGN FILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 1.320 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 1.320 5.440 ;
        END
    END VDD
END FILL2

MACRO FILL16
    CLASS CORE ;
    FOREIGN FILL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 10.560 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 10.560 5.440 ;
        END
    END VDD
END FILL16

MACRO FILL1
    CLASS CORE ;
    FOREIGN FILL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.660 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 0.660 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 0.660 5.440 ;
        END
    END VDD
END FILL1

MACRO RF2R1WX2
    CLASS CORE ;
    FOREIGN RF2R1WX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN WW
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 3.755 2.720 4.295 ;
        RECT  2.350 3.755 2.500 4.340 ;
        RECT  2.120 3.490 2.350 4.340 ;
        RECT  1.870 3.490 2.120 3.720 ;
        RECT  1.870 1.885 2.075 2.225 ;
        RECT  1.735 1.885 1.870 3.720 ;
        RECT  1.640 1.935 1.735 3.720 ;
        RECT  1.460 1.935 1.640 2.405 ;
        RECT  0.970 1.935 1.460 2.165 ;
        RECT  0.630 1.880 0.970 2.220 ;
        END
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.580 0.630 1.690 0.860 ;
        RECT  1.350 0.630 1.580 1.490 ;
        RECT  1.105 1.260 1.350 1.490 ;
        RECT  0.875 1.260 1.105 1.515 ;
        END
    END WB
    PIN R2W
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.990 0.630 8.465 1.220 ;
        END
    END R2W
    PIN R2B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  8.915 0.760 9.145 3.830 ;
        RECT  8.695 0.760 8.915 1.285 ;
        RECT  8.720 2.965 8.915 3.830 ;
        RECT  8.695 3.470 8.720 3.830 ;
        END
    END R2B
    PIN R1W
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 0.630 7.120 0.980 ;
        END
    END R1W
    PIN R1B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  6.150 0.865 6.260 1.675 ;
        RECT  6.150 2.770 6.260 3.580 ;
        RECT  5.920 0.865 6.150 3.580 ;
        RECT  5.725 0.865 5.920 1.540 ;
        RECT  5.495 1.260 5.725 1.540 ;
        END
    END R1B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.355 -0.400 10.560 0.400 ;
        RECT  10.015 -0.400 10.355 1.570 ;
        RECT  7.760 -0.400 10.015 0.400 ;
        RECT  7.420 -0.400 7.760 0.630 ;
        RECT  4.940 -0.400 7.420 0.400 ;
        RECT  4.600 -0.400 4.940 0.630 ;
        RECT  3.640 -0.400 4.600 0.400 ;
        RECT  3.300 -0.400 3.640 1.065 ;
        RECT  1.120 -0.400 3.300 0.400 ;
        RECT  0.780 -0.400 1.120 0.630 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.380 4.640 10.560 5.440 ;
        RECT  10.040 3.000 10.380 5.440 ;
        RECT  7.760 4.640 10.040 5.440 ;
        RECT  7.420 3.930 7.760 5.440 ;
        RECT  4.940 4.640 7.420 5.440 ;
        RECT  4.600 3.930 4.940 5.440 ;
        RECT  3.680 4.640 4.600 5.440 ;
        RECT  3.320 4.465 3.680 5.440 ;
        RECT  1.220 4.640 3.320 5.440 ;
        RECT  0.880 4.410 1.220 5.440 ;
        RECT  0.000 4.640 0.880 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.810 2.100 9.945 2.440 ;
        RECT  9.580 2.100 9.810 4.290 ;
        RECT  8.280 4.060 9.580 4.290 ;
        RECT  8.495 2.210 8.685 2.550 ;
        RECT  8.490 1.460 8.495 2.550 ;
        RECT  8.260 1.460 8.490 3.110 ;
        RECT  8.050 3.470 8.280 4.290 ;
        RECT  8.155 1.460 8.260 1.800 ;
        RECT  8.150 2.750 8.260 3.110 ;
        RECT  6.880 3.470 8.050 3.700 ;
        RECT  6.850 1.460 6.960 1.800 ;
        RECT  6.850 2.875 6.960 3.235 ;
        RECT  6.650 3.470 6.880 4.040 ;
        RECT  6.620 1.460 6.850 3.235 ;
        RECT  5.575 3.810 6.650 4.040 ;
        RECT  6.430 2.205 6.620 2.545 ;
        RECT  5.345 2.210 5.575 4.040 ;
        RECT  5.220 2.210 5.345 2.440 ;
        RECT  4.880 2.100 5.220 2.440 ;
        RECT  4.560 2.155 4.880 2.440 ;
        RECT  4.440 1.365 4.560 2.685 ;
        RECT  4.345 1.310 4.440 2.685 ;
        RECT  4.345 3.050 4.400 3.410 ;
        RECT  4.330 1.310 4.345 3.410 ;
        RECT  4.100 1.310 4.330 1.650 ;
        RECT  4.090 2.455 4.330 3.410 ;
        RECT  3.760 1.885 4.100 2.225 ;
        RECT  3.430 2.455 4.090 2.685 ;
        RECT  4.060 3.050 4.090 3.410 ;
        RECT  2.535 1.935 3.760 2.165 ;
        RECT  3.090 2.395 3.430 2.735 ;
        RECT  2.480 1.370 2.535 3.255 ;
        RECT  2.305 1.315 2.480 3.255 ;
        RECT  2.140 1.315 2.305 1.655 ;
        RECT  2.100 2.895 2.305 3.255 ;
        RECT  1.550 3.950 1.890 4.295 ;
        RECT  0.560 3.950 1.550 4.180 ;
        RECT  0.400 2.980 0.560 4.180 ;
        RECT  0.400 1.310 0.520 1.650 ;
        RECT  0.330 1.310 0.400 4.180 ;
        RECT  0.170 1.310 0.330 3.340 ;
    END
END RF2R1WX2

MACRO RF1R1WX2
    CLASS CORE ;
    FOREIGN RF1R1WX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN WW
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 3.480 2.735 4.000 ;
        RECT  2.425 3.480 2.505 3.780 ;
        RECT  1.745 3.480 2.425 3.710 ;
        RECT  1.840 1.610 2.015 2.610 ;
        RECT  1.785 1.610 1.840 2.660 ;
        RECT  1.745 2.380 1.785 2.660 ;
        RECT  1.515 2.380 1.745 3.710 ;
        RECT  1.460 2.380 1.515 2.660 ;
        RECT  0.825 2.405 1.460 2.635 ;
        RECT  0.595 2.405 0.825 2.775 ;
        END
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.965 1.285 1.195 2.105 ;
        RECT  0.875 1.285 0.965 1.515 ;
        END
    END WB
    PIN RWN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 3.500 6.460 3.780 ;
        RECT  6.080 3.500 6.310 4.235 ;
        RECT  4.835 4.005 6.080 4.235 ;
        RECT  4.390 4.005 4.835 4.370 ;
        END
    END RWN
    PIN RW
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 0.670 4.590 1.010 ;
        RECT  3.815 0.640 4.480 1.010 ;
        END
    END RW
    PIN RB
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.085 2.920 5.100 3.280 ;
        RECT  4.855 0.765 5.085 3.280 ;
        RECT  4.835 1.285 4.855 1.515 ;
        RECT  4.760 2.920 4.855 3.280 ;
        END
    END RB
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 -0.400 6.600 0.400 ;
        RECT  6.080 -0.400 6.420 1.585 ;
        RECT  3.585 -0.400 6.080 0.400 ;
        RECT  3.245 -0.400 3.585 1.030 ;
        RECT  1.320 -0.400 3.245 0.400 ;
        RECT  0.980 -0.400 1.320 0.645 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 4.640 6.600 5.440 ;
        RECT  6.080 4.465 6.420 5.440 ;
        RECT  3.485 4.640 6.080 5.440 ;
        RECT  3.145 3.700 3.485 5.440 ;
        RECT  1.280 4.640 3.145 5.440 ;
        RECT  0.940 4.400 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.790 2.100 6.050 2.440 ;
        RECT  5.710 2.100 5.790 3.740 ;
        RECT  5.560 2.205 5.710 3.740 ;
        RECT  4.340 3.510 5.560 3.740 ;
        RECT  4.285 1.340 4.500 2.880 ;
        RECT  4.285 3.250 4.340 3.740 ;
        RECT  4.270 1.340 4.285 3.740 ;
        RECT  4.065 1.340 4.270 1.680 ;
        RECT  4.055 2.650 4.270 3.740 ;
        RECT  3.370 2.650 4.055 2.880 ;
        RECT  4.000 3.250 4.055 3.610 ;
        RECT  3.700 1.910 4.040 2.250 ;
        RECT  2.475 1.960 3.700 2.190 ;
        RECT  3.030 2.540 3.370 2.880 ;
        RECT  2.475 0.970 2.480 1.310 ;
        RECT  2.245 0.970 2.475 3.250 ;
        RECT  2.140 0.970 2.245 1.310 ;
        RECT  2.060 3.020 2.245 3.250 ;
        RECT  1.745 4.085 2.120 4.315 ;
        RECT  1.515 3.940 1.745 4.315 ;
        RECT  0.465 3.940 1.515 4.170 ;
        RECT  0.365 0.870 0.520 1.100 ;
        RECT  0.365 3.170 0.465 4.170 ;
        RECT  0.235 0.870 0.365 4.170 ;
        RECT  0.135 0.870 0.235 3.400 ;
    END
END RF1R1WX2

MACRO XOR2XL
    CLASS CORE ;
    FOREIGN XOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 1.170 5.100 3.340 ;
        RECT  4.760 1.170 4.870 1.510 ;
        RECT  4.835 2.405 4.870 2.635 ;
        RECT  4.760 3.000 4.870 3.340 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 2.395 1.430 2.625 ;
        RECT  1.090 2.395 1.320 3.195 ;
        RECT  0.875 2.965 1.090 3.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 2.340 2.045 2.680 ;
        RECT  1.660 1.845 1.890 2.680 ;
        RECT  1.535 1.845 1.660 2.085 ;
        RECT  0.875 1.855 1.535 2.085 ;
        RECT  0.840 1.820 0.875 2.085 ;
        RECT  0.610 1.630 0.840 2.085 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 -0.400 5.280 0.400 ;
        RECT  4.200 -0.400 4.540 0.575 ;
        RECT  1.225 -0.400 4.200 0.400 ;
        RECT  0.885 -0.400 1.225 0.575 ;
        RECT  0.000 -0.400 0.885 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 4.640 5.280 5.440 ;
        RECT  4.200 4.465 4.540 5.440 ;
        RECT  1.150 4.640 4.200 5.440 ;
        RECT  0.810 4.465 1.150 5.440 ;
        RECT  0.000 4.640 0.810 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.475 1.740 4.635 2.080 ;
        RECT  4.245 0.815 4.475 2.080 ;
        RECT  2.965 0.815 4.245 1.045 ;
        RECT  3.670 3.605 4.010 4.160 ;
        RECT  3.675 1.275 3.905 3.315 ;
        RECT  3.400 1.275 3.675 1.505 ;
        RECT  3.455 2.950 3.675 3.315 ;
        RECT  2.505 3.605 3.670 3.835 ;
        RECT  1.610 4.090 3.300 4.320 ;
        RECT  2.735 0.815 2.965 3.370 ;
        RECT  1.685 0.630 2.505 0.860 ;
        RECT  2.275 1.305 2.505 3.835 ;
        RECT  1.800 1.305 2.275 1.535 ;
        RECT  1.800 3.130 2.275 3.470 ;
        RECT  1.455 0.630 1.685 1.035 ;
        RECT  1.380 3.790 1.610 4.320 ;
        RECT  0.520 0.805 1.455 1.035 ;
        RECT  0.520 3.790 1.380 4.020 ;
        RECT  0.380 0.805 0.520 1.345 ;
        RECT  0.380 3.400 0.520 4.020 ;
        RECT  0.290 0.805 0.380 4.020 ;
        RECT  0.150 1.115 0.290 3.785 ;
    END
END XOR2XL

MACRO XOR2X4
    CLASS CORE ;
    FOREIGN XOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR2XL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.190 1.410 10.420 4.340 ;
        RECT  10.020 1.410 10.190 1.750 ;
        RECT  10.040 2.940 10.190 4.340 ;
        RECT  10.020 3.050 10.040 3.525 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.100 1.490 2.440 ;
        RECT  0.875 2.100 1.105 2.635 ;
        RECT  0.550 2.100 0.875 2.440 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.475 2.310 7.705 2.635 ;
        RECT  7.060 2.310 7.475 2.540 ;
        RECT  6.720 2.200 7.060 2.540 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.220 0.400 ;
        RECT  10.700 -0.400 11.040 0.575 ;
        RECT  9.680 -0.400 10.700 0.400 ;
        RECT  9.340 -0.400 9.680 0.575 ;
        RECT  8.180 -0.400 9.340 0.400 ;
        RECT  7.840 -0.400 8.180 0.575 ;
        RECT  3.120 -0.400 7.840 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  1.800 -0.400 2.780 0.400 ;
        RECT  1.460 -0.400 1.800 1.020 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 1.020 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 4.640 11.220 5.440 ;
        RECT  10.700 4.465 11.040 5.440 ;
        RECT  9.680 4.640 10.700 5.440 ;
        RECT  9.340 4.465 9.680 5.440 ;
        RECT  8.240 4.640 9.340 5.440 ;
        RECT  7.900 4.465 8.240 5.440 ;
        RECT  3.120 4.640 7.900 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  1.800 4.640 2.780 5.440 ;
        RECT  1.460 4.090 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 4.090 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.755 2.210 9.960 2.550 ;
        RECT  9.525 0.865 9.755 2.550 ;
        RECT  7.460 0.865 9.525 1.095 ;
        RECT  8.770 1.410 9.000 3.380 ;
        RECT  8.660 1.410 8.770 1.885 ;
        RECT  8.660 3.040 8.770 3.380 ;
        RECT  6.740 1.655 8.660 1.885 ;
        RECT  8.415 2.330 8.540 2.670 ;
        RECT  8.185 2.330 8.415 4.185 ;
        RECT  6.740 3.955 8.185 4.185 ;
        RECT  7.120 0.865 7.460 1.250 ;
        RECT  7.120 3.280 7.460 3.620 ;
        RECT  6.020 0.865 7.120 1.095 ;
        RECT  6.085 3.340 7.120 3.570 ;
        RECT  6.405 1.340 6.740 1.885 ;
        RECT  6.400 3.800 6.740 4.185 ;
        RECT  6.400 1.340 6.405 3.070 ;
        RECT  6.175 1.655 6.400 3.070 ;
        RECT  3.525 3.955 6.400 4.185 ;
        RECT  5.300 2.840 6.175 3.070 ;
        RECT  5.680 3.340 6.085 3.725 ;
        RECT  5.885 0.865 6.020 1.330 ;
        RECT  5.655 0.865 5.885 1.825 ;
        RECT  4.645 3.495 5.680 3.725 ;
        RECT  4.645 1.595 5.655 1.825 ;
        RECT  4.960 0.865 5.300 1.280 ;
        RECT  4.960 2.840 5.300 3.180 ;
        RECT  2.440 0.865 4.960 1.095 ;
        RECT  4.580 1.595 4.645 3.725 ;
        RECT  4.415 1.455 4.580 3.725 ;
        RECT  4.230 1.455 4.415 1.825 ;
        RECT  4.240 3.350 4.415 3.725 ;
        RECT  3.825 2.155 4.125 2.555 ;
        RECT  3.825 1.420 3.880 1.760 ;
        RECT  3.825 3.000 3.880 3.340 ;
        RECT  3.595 1.420 3.825 3.340 ;
        RECT  3.540 1.420 3.595 1.760 ;
        RECT  3.540 3.000 3.595 3.340 ;
        RECT  3.295 3.570 3.525 4.185 ;
        RECT  2.440 3.570 3.295 3.800 ;
        RECT  2.210 0.865 2.440 3.800 ;
        RECT  2.100 1.420 2.210 1.760 ;
        RECT  2.100 3.040 2.210 3.380 ;
        RECT  1.160 1.420 2.100 1.650 ;
        RECT  1.160 3.150 2.100 3.380 ;
        RECT  0.820 1.420 1.160 1.760 ;
        RECT  0.820 3.040 1.160 3.380 ;
    END
END XOR2X4

MACRO XOR2X2
    CLASS CORE ;
    FOREIGN XOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR2XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.180 0.720 6.410 4.190 ;
        RECT  6.070 0.720 6.180 1.660 ;
        RECT  6.070 2.910 6.180 4.190 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 2.370 1.690 2.915 ;
        RECT  1.195 2.685 1.350 2.915 ;
        RECT  0.965 2.685 1.195 3.205 ;
        RECT  0.875 2.965 0.965 3.205 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.185 2.095 3.415 2.455 ;
        RECT  2.515 2.225 3.185 2.455 ;
        RECT  2.335 2.225 2.515 2.645 ;
        RECT  2.105 1.905 2.335 2.645 ;
        RECT  0.840 1.905 2.105 2.135 ;
        RECT  0.610 1.905 0.840 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.620 -0.400 6.600 0.400 ;
        RECT  5.280 -0.400 5.620 0.575 ;
        RECT  2.640 -0.400 5.280 0.400 ;
        RECT  2.300 -0.400 2.640 0.575 ;
        RECT  1.120 -0.400 2.300 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.610 4.640 6.600 5.440 ;
        RECT  5.270 4.465 5.610 5.440 ;
        RECT  2.560 4.640 5.270 5.440 ;
        RECT  2.220 3.740 2.560 5.440 ;
        RECT  1.120 4.640 2.220 5.440 ;
        RECT  0.780 3.740 1.120 5.440 ;
        RECT  0.000 4.640 0.780 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.805 1.985 5.945 2.345 ;
        RECT  5.575 0.890 5.805 2.345 ;
        RECT  4.335 0.890 5.575 1.120 ;
        RECT  5.045 2.185 5.275 4.175 ;
        RECT  3.280 3.945 5.045 4.175 ;
        RECT  4.565 1.410 4.795 3.370 ;
        RECT  4.105 0.890 4.335 3.520 ;
        RECT  3.720 0.890 4.105 1.230 ;
        RECT  4.000 3.290 4.105 3.520 ;
        RECT  3.660 3.290 4.000 3.630 ;
        RECT  3.645 1.545 3.875 2.975 ;
        RECT  3.470 1.545 3.645 1.775 ;
        RECT  3.280 2.745 3.645 2.975 ;
        RECT  3.340 0.865 3.470 1.775 ;
        RECT  3.240 0.685 3.340 1.775 ;
        RECT  3.050 2.745 3.280 4.175 ;
        RECT  3.000 0.685 3.240 1.095 ;
        RECT  2.940 3.010 3.050 3.950 ;
        RECT  1.880 0.865 3.000 1.095 ;
        RECT  2.630 1.340 2.970 1.680 ;
        RECT  1.840 3.215 2.940 3.445 ;
        RECT  0.520 1.395 2.630 1.625 ;
        RECT  1.540 0.810 1.880 1.150 ;
        RECT  1.610 3.215 1.840 3.800 ;
        RECT  1.500 3.460 1.610 3.800 ;
        RECT  0.380 1.180 0.520 1.625 ;
        RECT  0.380 2.870 0.520 3.210 ;
        RECT  0.380 3.990 0.505 4.330 ;
        RECT  0.150 1.180 0.380 4.330 ;
    END
END XOR2X2

MACRO XOR2X1
    CLASS CORE ;
    FOREIGN XOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 1.170 5.100 3.310 ;
        RECT  4.760 1.170 4.870 1.510 ;
        RECT  4.835 2.405 4.870 3.310 ;
        RECT  4.760 2.970 4.835 3.310 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 2.395 1.430 2.625 ;
        RECT  1.090 2.395 1.320 3.195 ;
        RECT  0.875 2.965 1.090 3.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 2.340 2.045 2.680 ;
        RECT  1.660 1.845 1.890 2.680 ;
        RECT  1.535 1.845 1.660 2.085 ;
        RECT  0.875 1.855 1.535 2.085 ;
        RECT  0.840 1.820 0.875 2.085 ;
        RECT  0.610 1.630 0.840 2.085 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 -0.400 5.280 0.400 ;
        RECT  4.200 -0.400 4.540 0.575 ;
        RECT  1.225 -0.400 4.200 0.400 ;
        RECT  0.885 -0.400 1.225 0.575 ;
        RECT  0.000 -0.400 0.885 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 4.640 5.280 5.440 ;
        RECT  4.200 4.465 4.540 5.440 ;
        RECT  1.150 4.640 4.200 5.440 ;
        RECT  0.810 4.465 1.150 5.440 ;
        RECT  0.000 4.640 0.810 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.475 1.790 4.635 2.130 ;
        RECT  4.245 0.815 4.475 2.130 ;
        RECT  3.005 0.815 4.245 1.045 ;
        RECT  3.670 3.605 4.010 4.090 ;
        RECT  3.675 1.275 3.905 3.315 ;
        RECT  3.440 1.275 3.675 1.505 ;
        RECT  3.495 2.950 3.675 3.315 ;
        RECT  2.505 3.605 3.670 3.835 ;
        RECT  1.610 4.090 3.300 4.320 ;
        RECT  2.775 0.815 3.005 3.370 ;
        RECT  1.685 0.630 2.545 0.860 ;
        RECT  2.275 1.305 2.505 3.835 ;
        RECT  1.800 1.305 2.275 1.535 ;
        RECT  1.800 3.130 2.275 3.470 ;
        RECT  1.455 0.630 1.685 1.035 ;
        RECT  1.380 3.790 1.610 4.320 ;
        RECT  0.520 0.805 1.455 1.035 ;
        RECT  0.520 3.790 1.380 4.020 ;
        RECT  0.380 0.805 0.520 1.315 ;
        RECT  0.380 3.400 0.520 4.020 ;
        RECT  0.290 0.805 0.380 4.020 ;
        RECT  0.150 1.085 0.290 3.785 ;
    END
END XOR2X1

MACRO XNOR2XL
    CLASS CORE ;
    FOREIGN XNOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 1.150 5.100 3.320 ;
        RECT  4.760 1.150 4.870 1.490 ;
        RECT  4.835 2.405 4.870 3.320 ;
        RECT  4.815 2.975 4.835 3.320 ;
        RECT  4.760 2.980 4.815 3.320 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 2.395 1.430 2.625 ;
        RECT  1.090 2.395 1.320 3.195 ;
        RECT  0.875 2.965 1.090 3.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 2.180 2.045 2.540 ;
        RECT  1.660 1.845 1.890 2.540 ;
        RECT  1.535 1.845 1.660 2.085 ;
        RECT  0.875 1.855 1.535 2.085 ;
        RECT  0.840 1.820 0.875 2.085 ;
        RECT  0.610 1.630 0.840 2.085 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 -0.400 5.280 0.400 ;
        RECT  4.200 -0.400 4.540 0.575 ;
        RECT  1.225 -0.400 4.200 0.400 ;
        RECT  0.885 -0.400 1.225 0.575 ;
        RECT  0.000 -0.400 0.885 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 4.640 5.280 5.440 ;
        RECT  4.200 4.465 4.540 5.440 ;
        RECT  1.150 4.640 4.200 5.440 ;
        RECT  0.810 4.465 1.150 5.440 ;
        RECT  0.000 4.640 0.810 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.530 1.790 4.635 2.130 ;
        RECT  4.300 1.790 4.530 3.775 ;
        RECT  2.965 3.545 4.300 3.775 ;
        RECT  2.505 4.005 4.010 4.235 ;
        RECT  3.675 1.240 3.905 3.265 ;
        RECT  3.400 1.240 3.675 1.580 ;
        RECT  3.440 3.035 3.675 3.265 ;
        RECT  1.685 0.645 3.260 0.875 ;
        RECT  2.735 1.225 2.965 3.775 ;
        RECT  2.275 1.295 2.505 4.235 ;
        RECT  1.800 1.295 2.275 1.525 ;
        RECT  1.800 3.130 2.275 3.470 ;
        RECT  1.815 3.790 2.045 4.270 ;
        RECT  0.520 3.790 1.815 4.020 ;
        RECT  1.455 0.645 1.685 1.035 ;
        RECT  0.520 0.805 1.455 1.035 ;
        RECT  0.380 0.805 0.520 1.400 ;
        RECT  0.380 3.400 0.520 4.020 ;
        RECT  0.290 0.805 0.380 4.020 ;
        RECT  0.150 1.060 0.290 3.785 ;
    END
END XNOR2XL

MACRO XNOR2X4
    CLASS CORE ;
    FOREIGN XNOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR2XL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.190 1.410 10.420 4.340 ;
        RECT  10.020 1.410 10.190 1.750 ;
        RECT  10.040 2.940 10.190 4.340 ;
        RECT  10.020 3.050 10.040 3.390 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.100 1.490 2.440 ;
        RECT  0.875 2.100 1.105 2.635 ;
        RECT  0.550 2.100 0.875 2.440 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.205 2.170 3.540 2.510 ;
        RECT  2.855 2.170 3.205 2.635 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.220 0.400 ;
        RECT  10.700 -0.400 11.040 0.575 ;
        RECT  9.680 -0.400 10.700 0.400 ;
        RECT  9.340 -0.400 9.680 0.575 ;
        RECT  8.180 -0.400 9.340 0.400 ;
        RECT  7.840 -0.400 8.180 0.575 ;
        RECT  3.120 -0.400 7.840 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  1.800 -0.400 2.780 0.400 ;
        RECT  1.460 -0.400 1.800 1.020 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 1.020 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 4.640 11.220 5.440 ;
        RECT  10.700 4.465 11.040 5.440 ;
        RECT  9.680 4.640 10.700 5.440 ;
        RECT  9.340 4.465 9.680 5.440 ;
        RECT  8.240 4.640 9.340 5.440 ;
        RECT  7.900 4.465 8.240 5.440 ;
        RECT  3.120 4.640 7.900 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  1.800 4.640 2.780 5.440 ;
        RECT  1.460 4.090 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 4.090 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.755 2.210 9.960 2.550 ;
        RECT  9.525 0.865 9.755 4.035 ;
        RECT  7.460 0.865 9.525 1.095 ;
        RECT  4.240 3.805 9.525 4.035 ;
        RECT  8.770 1.410 9.000 3.380 ;
        RECT  8.660 1.410 8.770 1.885 ;
        RECT  8.660 3.040 8.770 3.380 ;
        RECT  7.620 1.655 8.660 1.885 ;
        RECT  8.415 2.330 8.540 2.670 ;
        RECT  8.185 2.330 8.415 3.575 ;
        RECT  2.440 3.345 8.185 3.575 ;
        RECT  7.390 1.655 7.620 3.005 ;
        RECT  7.120 0.865 7.460 1.250 ;
        RECT  6.740 1.655 7.390 1.885 ;
        RECT  5.300 2.775 7.390 3.005 ;
        RECT  6.020 0.865 7.120 1.095 ;
        RECT  6.720 2.200 7.060 2.540 ;
        RECT  6.445 1.340 6.740 1.885 ;
        RECT  4.000 2.255 6.720 2.485 ;
        RECT  6.400 1.340 6.445 1.680 ;
        RECT  5.885 0.865 6.020 1.330 ;
        RECT  5.655 0.865 5.885 1.685 ;
        RECT  4.240 1.455 5.655 1.685 ;
        RECT  4.960 0.865 5.300 1.225 ;
        RECT  4.960 2.775 5.300 3.115 ;
        RECT  2.440 0.865 4.960 1.095 ;
        RECT  3.770 1.420 4.000 3.080 ;
        RECT  3.540 1.420 3.770 1.760 ;
        RECT  3.540 2.740 3.770 3.080 ;
        RECT  2.210 0.865 2.440 3.575 ;
        RECT  2.100 1.420 2.210 1.760 ;
        RECT  2.100 3.040 2.210 3.380 ;
        RECT  1.160 1.420 2.100 1.650 ;
        RECT  1.160 3.150 2.100 3.380 ;
        RECT  0.820 1.420 1.160 1.760 ;
        RECT  0.820 3.040 1.160 3.380 ;
    END
END XNOR2X4

MACRO XNOR2X2
    CLASS CORE ;
    FOREIGN XNOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR2XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.070 0.720 7.080 1.660 ;
        RECT  6.840 0.720 7.070 4.190 ;
        RECT  6.740 0.720 6.840 1.660 ;
        RECT  6.730 2.910 6.840 4.190 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 2.370 1.890 2.710 ;
        RECT  1.550 2.370 1.780 2.915 ;
        RECT  1.460 2.635 1.550 2.915 ;
        RECT  1.195 2.685 1.460 2.915 ;
        RECT  0.965 2.685 1.195 3.205 ;
        RECT  0.875 2.965 0.965 3.205 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.845 1.965 4.075 2.455 ;
        RECT  3.175 2.225 3.845 2.455 ;
        RECT  2.945 2.225 3.175 2.645 ;
        RECT  2.425 2.415 2.945 2.645 ;
        RECT  2.350 2.405 2.425 2.645 ;
        RECT  2.120 1.905 2.350 2.645 ;
        RECT  0.840 1.905 2.120 2.135 ;
        RECT  0.610 1.905 0.840 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 -0.400 7.260 0.400 ;
        RECT  5.980 -0.400 6.320 0.575 ;
        RECT  2.940 -0.400 5.980 0.400 ;
        RECT  2.600 -0.400 2.940 0.575 ;
        RECT  1.400 -0.400 2.600 0.400 ;
        RECT  1.060 -0.400 1.400 0.575 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.270 4.640 7.260 5.440 ;
        RECT  5.930 4.465 6.270 5.440 ;
        RECT  2.860 4.640 5.930 5.440 ;
        RECT  2.520 3.740 2.860 5.440 ;
        RECT  1.380 4.640 2.520 5.440 ;
        RECT  1.040 3.740 1.380 5.440 ;
        RECT  0.000 4.640 1.040 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.465 1.980 6.605 2.345 ;
        RECT  6.235 0.825 6.465 2.345 ;
        RECT  4.995 0.825 6.235 1.055 ;
        RECT  5.705 2.185 5.935 4.175 ;
        RECT  3.710 3.945 5.705 4.175 ;
        RECT  5.225 1.285 5.455 3.370 ;
        RECT  4.765 0.825 4.995 3.520 ;
        RECT  4.380 0.825 4.765 1.270 ;
        RECT  4.660 3.290 4.765 3.520 ;
        RECT  4.320 3.290 4.660 3.630 ;
        RECT  4.305 1.500 4.535 2.975 ;
        RECT  3.945 1.500 4.305 1.730 ;
        RECT  3.710 2.745 4.305 2.975 ;
        RECT  3.715 0.835 3.945 1.730 ;
        RECT  2.180 0.835 3.715 1.065 ;
        RECT  3.480 2.745 3.710 4.175 ;
        RECT  3.365 3.010 3.480 3.950 ;
        RECT  3.130 1.295 3.470 1.635 ;
        RECT  2.140 3.215 3.365 3.445 ;
        RECT  0.520 1.350 3.130 1.580 ;
        RECT  1.840 0.780 2.180 1.120 ;
        RECT  1.910 3.215 2.140 3.800 ;
        RECT  1.800 3.460 1.910 3.800 ;
        RECT  0.380 1.180 0.520 1.580 ;
        RECT  0.380 2.870 0.520 3.210 ;
        RECT  0.380 3.990 0.505 4.330 ;
        RECT  0.150 1.180 0.380 4.330 ;
    END
END XNOR2X2

MACRO XNOR2X1
    CLASS CORE ;
    FOREIGN XNOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 1.170 5.100 3.310 ;
        RECT  4.760 1.170 4.870 1.510 ;
        RECT  4.835 2.405 4.870 3.310 ;
        RECT  4.760 2.970 4.835 3.310 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 2.330 1.430 2.670 ;
        RECT  1.090 2.330 1.320 3.195 ;
        RECT  0.875 2.965 1.090 3.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 2.340 2.045 2.680 ;
        RECT  1.660 1.845 1.890 2.680 ;
        RECT  1.535 1.845 1.660 2.085 ;
        RECT  0.875 1.855 1.535 2.085 ;
        RECT  0.840 1.845 0.875 2.085 ;
        RECT  0.610 1.630 0.840 2.085 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 -0.400 5.280 0.400 ;
        RECT  4.200 -0.400 4.540 0.575 ;
        RECT  1.225 -0.400 4.200 0.400 ;
        RECT  0.885 -0.400 1.225 0.575 ;
        RECT  0.000 -0.400 0.885 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 4.640 5.280 5.440 ;
        RECT  4.200 4.465 4.540 5.440 ;
        RECT  1.200 4.640 4.200 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.530 1.790 4.635 2.130 ;
        RECT  4.300 1.790 4.530 3.490 ;
        RECT  2.965 3.260 4.300 3.490 ;
        RECT  3.670 3.720 4.010 4.090 ;
        RECT  3.675 1.240 3.905 3.025 ;
        RECT  3.495 1.240 3.675 1.580 ;
        RECT  3.440 2.795 3.675 3.025 ;
        RECT  2.505 3.720 3.670 3.950 ;
        RECT  2.920 0.665 3.260 1.005 ;
        RECT  2.735 1.240 2.965 3.490 ;
        RECT  1.685 0.775 2.920 1.005 ;
        RECT  1.945 4.180 2.710 4.410 ;
        RECT  2.275 1.350 2.505 3.950 ;
        RECT  2.140 1.350 2.275 1.580 ;
        RECT  1.800 3.130 2.275 3.470 ;
        RECT  1.800 1.240 2.140 1.580 ;
        RECT  1.715 3.790 1.945 4.410 ;
        RECT  0.520 3.790 1.715 4.020 ;
        RECT  1.455 0.775 1.685 1.035 ;
        RECT  0.520 0.805 1.455 1.035 ;
        RECT  0.380 0.805 0.520 1.370 ;
        RECT  0.380 3.400 0.520 4.020 ;
        RECT  0.290 0.805 0.380 4.020 ;
        RECT  0.150 0.805 0.290 3.785 ;
    END
END XNOR2X1

MACRO TLATSRXL
    CLASS CORE ;
    FOREIGN TLATSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.105 0.555 2.445 ;
        RECT  0.140 1.840 0.545 2.445 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.510 1.845 3.820 2.500 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.005 1.240 11.040 1.580 ;
        RECT  11.005 3.020 11.040 3.360 ;
        RECT  10.775 1.240 11.005 3.360 ;
        RECT  10.700 1.240 10.775 1.580 ;
        RECT  10.700 3.020 10.775 3.360 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.640 2.965 9.685 3.205 ;
        RECT  9.620 2.965 9.640 3.310 ;
        RECT  9.390 1.430 9.620 3.310 ;
        RECT  9.280 1.430 9.390 1.770 ;
        RECT  9.300 2.970 9.390 3.310 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.600 1.930 6.940 2.270 ;
        RECT  6.385 1.930 6.600 2.160 ;
        RECT  6.155 1.845 6.385 2.160 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.900 3.085 2.660 ;
        RECT  2.580 1.900 2.780 2.240 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 -0.400 11.220 0.400 ;
        RECT  9.980 -0.400 10.320 0.575 ;
        RECT  8.820 -0.400 9.980 0.400 ;
        RECT  8.480 -0.400 8.820 0.575 ;
        RECT  6.320 -0.400 8.480 0.400 ;
        RECT  5.980 -0.400 6.320 0.575 ;
        RECT  2.720 -0.400 5.980 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  0.520 -0.400 2.380 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.385 4.640 11.220 5.440 ;
        RECT  9.975 4.465 10.385 5.440 ;
        RECT  8.880 4.640 9.975 5.440 ;
        RECT  8.540 4.465 8.880 5.440 ;
        RECT  6.860 4.640 8.540 5.440 ;
        RECT  6.520 4.465 6.860 5.440 ;
        RECT  3.500 4.640 6.520 5.440 ;
        RECT  3.160 4.135 3.500 5.440 ;
        RECT  0.520 4.640 3.160 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.185 0.805 10.415 4.015 ;
        RECT  9.620 0.805 10.185 1.035 ;
        RECT  9.640 3.785 10.185 4.015 ;
        RECT  9.410 3.785 9.640 4.365 ;
        RECT  9.280 0.665 9.620 1.035 ;
        RECT  9.300 4.005 9.410 4.365 ;
        RECT  5.990 4.005 9.300 4.235 ;
        RECT  9.025 2.090 9.160 2.430 ;
        RECT  8.795 2.090 9.025 3.775 ;
        RECT  4.860 3.545 8.795 3.775 ;
        RECT  7.965 0.745 8.195 3.270 ;
        RECT  7.680 0.745 7.965 1.085 ;
        RECT  7.820 2.930 7.965 3.270 ;
        RECT  7.485 1.900 7.730 2.240 ;
        RECT  5.655 0.855 7.680 1.085 ;
        RECT  7.255 1.315 7.485 3.315 ;
        RECT  6.980 1.315 7.255 1.545 ;
        RECT  5.585 3.085 7.255 3.315 ;
        RECT  5.425 0.855 5.655 2.665 ;
        RECT  5.355 2.895 5.585 3.315 ;
        RECT  4.850 2.435 5.425 2.665 ;
        RECT  4.305 2.895 5.355 3.125 ;
        RECT  4.670 1.710 5.010 2.050 ;
        RECT  4.520 3.365 4.860 3.775 ;
        RECT  4.305 1.765 4.670 2.050 ;
        RECT  4.260 1.130 4.600 1.470 ;
        RECT  1.820 3.545 4.520 3.775 ;
        RECT  4.075 1.765 4.305 3.125 ;
        RECT  2.595 1.240 4.260 1.470 ;
        RECT  2.475 2.895 4.075 3.125 ;
        RECT  2.365 1.240 2.595 1.545 ;
        RECT  2.245 2.470 2.475 3.125 ;
        RECT  1.620 1.315 2.365 1.545 ;
        RECT  2.190 2.470 2.245 2.700 ;
        RECT  1.850 2.360 2.190 2.700 ;
        RECT  1.620 0.730 1.960 1.070 ;
        RECT  1.620 3.110 1.820 3.775 ;
        RECT  1.290 4.020 1.630 4.360 ;
        RECT  1.120 0.840 1.620 1.070 ;
        RECT  1.590 1.315 1.620 3.775 ;
        RECT  1.390 1.315 1.590 3.450 ;
        RECT  1.120 4.020 1.290 4.250 ;
        RECT  0.890 0.840 1.120 4.250 ;
        RECT  0.780 1.290 0.890 1.630 ;
        RECT  0.780 3.000 0.890 3.340 ;
    END
END TLATSRXL

MACRO TLATSRX4
    CLASS CORE ;
    FOREIGN TLATSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.790 1.900 1.105 2.635 ;
        RECT  0.710 1.900 0.790 2.405 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.760 1.765 9.100 2.395 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.680 1.820 15.700 3.220 ;
        RECT  15.340 1.260 15.680 3.220 ;
        RECT  15.320 1.820 15.340 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.380 1.260 14.400 1.600 ;
        RECT  14.380 2.880 14.400 3.220 ;
        RECT  14.060 1.260 14.380 3.220 ;
        RECT  14.000 1.820 14.060 3.220 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  10.080 1.845 10.420 2.505 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.950 2.295 5.290 2.635 ;
        RECT  3.745 2.350 4.950 2.580 ;
        RECT  3.515 1.845 3.745 2.580 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 -0.400 16.500 0.400 ;
        RECT  15.980 -0.400 16.320 0.950 ;
        RECT  15.040 -0.400 15.980 0.400 ;
        RECT  14.700 -0.400 15.040 0.950 ;
        RECT  13.720 -0.400 14.700 0.400 ;
        RECT  13.380 -0.400 13.720 0.575 ;
        RECT  12.220 -0.400 13.380 0.400 ;
        RECT  11.880 -0.400 12.220 0.575 ;
        RECT  9.940 -0.400 11.880 0.400 ;
        RECT  9.600 -0.400 9.940 0.575 ;
        RECT  6.100 -0.400 9.600 0.400 ;
        RECT  5.760 -0.400 6.100 0.920 ;
        RECT  2.965 -0.400 5.760 0.400 ;
        RECT  2.625 -0.400 2.965 0.575 ;
        RECT  1.280 -0.400 2.625 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 4.640 16.500 5.440 ;
        RECT  15.980 4.090 16.320 5.440 ;
        RECT  15.040 4.640 15.980 5.440 ;
        RECT  14.700 4.090 15.040 5.440 ;
        RECT  13.720 4.640 14.700 5.440 ;
        RECT  13.380 4.465 13.720 5.440 ;
        RECT  12.200 4.640 13.380 5.440 ;
        RECT  11.860 4.465 12.200 5.440 ;
        RECT  10.340 4.640 11.860 5.440 ;
        RECT  10.000 4.465 10.340 5.440 ;
        RECT  6.980 4.640 10.000 5.440 ;
        RECT  6.640 4.465 6.980 5.440 ;
        RECT  1.200 4.640 6.640 5.440 ;
        RECT  0.860 3.850 1.200 5.440 ;
        RECT  0.820 3.850 0.860 4.190 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.160 2.070 16.270 2.410 ;
        RECT  15.930 2.070 16.160 3.785 ;
        RECT  12.905 3.555 15.930 3.785 ;
        RECT  13.465 1.370 13.695 3.015 ;
        RECT  12.980 1.370 13.465 1.600 ;
        RECT  12.905 2.785 13.465 3.015 ;
        RECT  12.395 2.080 13.190 2.420 ;
        RECT  12.640 1.260 12.980 1.600 ;
        RECT  12.675 2.785 12.905 4.225 ;
        RECT  9.470 3.995 12.675 4.225 ;
        RECT  12.165 2.080 12.395 3.655 ;
        RECT  2.545 3.425 12.165 3.655 ;
        RECT  11.645 1.215 11.875 3.085 ;
        RECT  11.460 1.215 11.645 1.445 ;
        RECT  11.640 2.855 11.645 3.085 ;
        RECT  11.300 2.855 11.640 3.195 ;
        RECT  11.350 1.105 11.460 1.445 ;
        RECT  10.955 1.685 11.355 2.075 ;
        RECT  11.120 0.805 11.350 1.445 ;
        RECT  9.345 0.805 11.120 1.035 ;
        RECT  10.890 1.685 10.955 3.195 ;
        RECT  10.660 1.265 10.890 3.195 ;
        RECT  10.400 1.265 10.660 1.495 ;
        RECT  8.375 2.965 10.660 3.195 ;
        RECT  9.115 0.805 9.345 1.355 ;
        RECT  7.540 4.180 9.140 4.410 ;
        RECT  7.720 1.125 9.115 1.355 ;
        RECT  8.375 1.585 8.430 1.925 ;
        RECT  8.145 1.585 8.375 3.195 ;
        RECT  8.090 1.585 8.145 1.925 ;
        RECT  3.130 2.965 8.145 3.195 ;
        RECT  6.985 0.665 8.020 0.895 ;
        RECT  7.490 1.125 7.720 2.355 ;
        RECT  7.310 3.945 7.540 4.410 ;
        RECT  7.380 1.835 7.490 2.355 ;
        RECT  4.550 1.835 7.380 2.065 ;
        RECT  6.065 3.945 7.310 4.175 ;
        RECT  6.755 0.665 6.985 1.385 ;
        RECT  2.545 1.155 6.755 1.385 ;
        RECT  5.835 3.945 6.065 4.355 ;
        RECT  1.865 4.125 5.835 4.355 ;
        RECT  4.210 1.780 4.550 2.120 ;
        RECT  2.900 2.210 3.130 3.195 ;
        RECT  2.790 2.210 2.900 2.550 ;
        RECT  2.315 1.155 2.545 3.655 ;
        RECT  1.800 1.155 2.315 1.495 ;
        RECT  1.865 1.790 2.000 2.130 ;
        RECT  1.635 1.790 1.865 4.355 ;
        RECT  1.565 1.790 1.635 2.020 ;
        RECT  0.520 2.975 1.635 3.245 ;
        RECT  1.335 1.415 1.565 2.020 ;
        RECT  0.520 1.415 1.335 1.645 ;
        RECT  0.180 0.835 0.520 1.645 ;
        RECT  0.180 2.905 0.520 3.245 ;
    END
END TLATSRX4

MACRO TLATSRX2
    CLASS CORE ;
    FOREIGN TLATSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 2.170 0.560 2.510 ;
        RECT  0.215 1.845 0.550 2.510 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 1.845 4.405 2.100 ;
        RECT  3.705 1.845 3.990 2.330 ;
        RECT  3.650 1.990 3.705 2.330 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.360 0.805 11.700 4.115 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.260 2.965 10.345 3.195 ;
        RECT  10.180 2.635 10.260 3.195 ;
        RECT  9.975 1.360 10.180 3.195 ;
        RECT  9.950 1.360 9.975 3.180 ;
        RECT  9.840 1.360 9.950 1.700 ;
        RECT  9.920 2.840 9.950 3.180 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.655 2.320 6.930 2.660 ;
        RECT  6.425 1.845 6.655 2.660 ;
        RECT  6.155 1.845 6.425 2.075 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.980 1.845 3.320 2.445 ;
        RECT  2.855 1.845 2.980 2.075 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.940 -0.400 11.880 0.400 ;
        RECT  10.600 -0.400 10.940 0.575 ;
        RECT  8.820 -0.400 10.600 0.400 ;
        RECT  8.480 -0.400 8.820 0.575 ;
        RECT  6.780 -0.400 8.480 0.400 ;
        RECT  6.440 -0.400 6.780 0.575 ;
        RECT  2.830 -0.400 6.440 0.400 ;
        RECT  2.490 -0.400 2.830 0.575 ;
        RECT  0.520 -0.400 2.490 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.980 4.640 11.880 5.440 ;
        RECT  10.640 4.090 10.980 5.440 ;
        RECT  8.800 4.640 10.640 5.440 ;
        RECT  8.460 4.465 8.800 5.440 ;
        RECT  6.900 4.640 8.460 5.440 ;
        RECT  6.560 4.465 6.900 5.440 ;
        RECT  3.620 4.640 6.560 5.440 ;
        RECT  3.280 3.740 3.620 5.440 ;
        RECT  0.520 4.640 3.280 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.900 0.885 11.130 3.835 ;
        RECT  9.480 0.885 10.900 1.115 ;
        RECT  9.560 3.605 10.900 3.835 ;
        RECT  9.220 2.070 9.560 2.410 ;
        RECT  9.450 3.090 9.560 3.835 ;
        RECT  9.140 0.885 9.480 1.430 ;
        RECT  9.220 3.090 9.450 4.235 ;
        RECT  8.765 2.180 9.220 2.410 ;
        RECT  6.030 4.005 9.220 4.235 ;
        RECT  8.535 2.180 8.765 3.655 ;
        RECT  4.900 3.425 8.535 3.655 ;
        RECT  8.065 1.095 8.245 3.190 ;
        RECT  8.015 0.875 8.065 3.190 ;
        RECT  7.780 0.875 8.015 1.440 ;
        RECT  7.860 2.850 8.015 3.190 ;
        RECT  5.755 0.875 7.780 1.105 ;
        RECT  7.500 1.930 7.780 2.270 ;
        RECT  7.270 1.360 7.500 3.190 ;
        RECT  7.080 1.360 7.270 1.700 ;
        RECT  7.160 2.850 7.270 3.190 ;
        RECT  5.590 2.905 7.160 3.135 ;
        RECT  5.590 0.875 5.755 2.505 ;
        RECT  5.525 0.875 5.590 2.560 ;
        RECT  5.360 2.790 5.590 3.135 ;
        RECT  5.250 2.220 5.525 2.560 ;
        RECT  5.015 2.790 5.360 3.020 ;
        RECT  5.015 1.550 5.270 1.890 ;
        RECT  4.785 1.550 5.015 3.020 ;
        RECT  4.560 0.960 4.900 1.300 ;
        RECT  4.560 3.260 4.900 3.710 ;
        RECT  2.550 2.755 4.785 2.985 ;
        RECT  3.430 1.070 4.560 1.300 ;
        RECT  1.780 3.260 4.560 3.490 ;
        RECT  3.200 1.070 3.430 1.440 ;
        RECT  1.880 1.210 3.200 1.440 ;
        RECT  2.320 2.320 2.550 2.985 ;
        RECT  2.150 2.320 2.320 2.550 ;
        RECT  1.810 2.210 2.150 2.550 ;
        RECT  1.580 1.085 1.880 1.440 ;
        RECT  1.580 3.000 1.780 3.810 ;
        RECT  1.540 1.085 1.580 3.810 ;
        RECT  1.440 1.210 1.540 3.810 ;
        RECT  1.350 1.210 1.440 3.600 ;
        RECT  1.080 0.720 1.270 0.950 ;
        RECT  0.850 0.720 1.080 3.735 ;
        RECT  0.740 1.245 0.850 1.585 ;
        RECT  0.740 2.925 0.850 3.735 ;
    END
END TLATSRX2

MACRO TLATSRX1
    CLASS CORE ;
    FOREIGN TLATSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSRXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.105 0.555 2.445 ;
        RECT  0.140 1.840 0.545 2.445 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 2.130 3.850 2.470 ;
        RECT  3.510 1.845 3.820 2.470 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.005 1.310 11.040 1.845 ;
        RECT  11.005 3.020 11.040 3.360 ;
        RECT  10.775 1.310 11.005 3.360 ;
        RECT  10.700 1.310 10.775 1.820 ;
        RECT  10.700 3.020 10.775 3.360 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.640 2.965 9.685 3.205 ;
        RECT  9.620 2.965 9.640 3.310 ;
        RECT  9.390 1.430 9.620 3.310 ;
        RECT  9.280 1.430 9.390 1.770 ;
        RECT  9.300 2.970 9.390 3.310 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 1.930 6.900 2.270 ;
        RECT  6.385 1.930 6.560 2.160 ;
        RECT  6.155 1.845 6.385 2.160 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.900 3.085 2.660 ;
        RECT  2.580 1.900 2.780 2.240 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 -0.400 11.220 0.400 ;
        RECT  9.980 -0.400 10.320 0.575 ;
        RECT  8.820 -0.400 9.980 0.400 ;
        RECT  8.480 -0.400 8.820 0.575 ;
        RECT  6.320 -0.400 8.480 0.400 ;
        RECT  5.980 -0.400 6.320 0.575 ;
        RECT  2.720 -0.400 5.980 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  0.520 -0.400 2.380 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.395 4.640 11.220 5.440 ;
        RECT  9.980 4.465 10.395 5.440 ;
        RECT  8.880 4.640 9.980 5.440 ;
        RECT  8.540 4.465 8.880 5.440 ;
        RECT  6.820 4.640 8.540 5.440 ;
        RECT  6.480 4.465 6.820 5.440 ;
        RECT  3.500 4.640 6.480 5.440 ;
        RECT  3.160 4.135 3.500 5.440 ;
        RECT  0.520 4.640 3.160 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.185 0.805 10.415 4.235 ;
        RECT  9.620 0.805 10.185 1.035 ;
        RECT  9.640 4.005 10.185 4.235 ;
        RECT  9.300 4.005 9.640 4.365 ;
        RECT  9.280 0.635 9.620 1.035 ;
        RECT  5.950 4.005 9.300 4.235 ;
        RECT  9.025 2.090 9.160 2.430 ;
        RECT  8.795 2.090 9.025 3.775 ;
        RECT  4.820 3.545 8.795 3.775 ;
        RECT  7.965 0.765 8.195 3.170 ;
        RECT  7.680 0.765 7.965 1.105 ;
        RECT  7.780 2.830 7.965 3.170 ;
        RECT  7.485 1.900 7.730 2.240 ;
        RECT  5.655 0.875 7.680 1.105 ;
        RECT  7.255 1.365 7.485 3.315 ;
        RECT  6.880 1.365 7.255 1.595 ;
        RECT  5.585 3.085 7.255 3.315 ;
        RECT  5.425 0.875 5.655 2.665 ;
        RECT  5.355 2.910 5.585 3.315 ;
        RECT  4.850 2.435 5.425 2.665 ;
        RECT  4.450 2.910 5.355 3.140 ;
        RECT  4.670 1.710 5.010 2.050 ;
        RECT  4.480 3.370 4.820 3.775 ;
        RECT  4.450 1.820 4.670 2.050 ;
        RECT  4.260 1.040 4.600 1.380 ;
        RECT  1.820 3.545 4.480 3.775 ;
        RECT  4.220 1.820 4.450 3.140 ;
        RECT  2.595 1.150 4.260 1.380 ;
        RECT  2.475 2.905 4.220 3.135 ;
        RECT  2.365 1.150 2.595 1.545 ;
        RECT  2.245 2.470 2.475 3.135 ;
        RECT  1.620 1.315 2.365 1.545 ;
        RECT  2.190 2.470 2.245 2.700 ;
        RECT  1.850 2.360 2.190 2.700 ;
        RECT  1.620 0.730 1.960 1.070 ;
        RECT  1.620 3.110 1.820 3.775 ;
        RECT  1.290 4.020 1.630 4.360 ;
        RECT  1.120 0.840 1.620 1.070 ;
        RECT  1.590 1.315 1.620 3.775 ;
        RECT  1.390 1.315 1.590 3.450 ;
        RECT  1.120 4.020 1.290 4.250 ;
        RECT  0.890 0.840 1.120 4.250 ;
        RECT  0.780 1.290 0.890 1.630 ;
        RECT  0.780 2.930 0.890 3.270 ;
    END
END TLATSRX1

MACRO TLATSXL
    CLASS CORE ;
    FOREIGN TLATSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 2.015 0.560 2.355 ;
        RECT  0.140 1.820 0.550 2.355 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 1.270 10.360 1.845 ;
        RECT  10.345 3.020 10.360 3.360 ;
        RECT  10.115 1.270 10.345 3.360 ;
        RECT  10.040 1.270 10.115 1.820 ;
        RECT  10.020 3.020 10.115 3.360 ;
        RECT  10.020 1.270 10.040 1.610 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.925 1.400 9.155 3.310 ;
        RECT  8.640 1.400 8.925 1.740 ;
        RECT  8.680 2.940 8.925 3.310 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.890 1.500 6.230 1.840 ;
        RECT  5.725 1.500 5.890 1.730 ;
        RECT  5.495 1.285 5.725 1.730 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.710 1.805 3.310 2.185 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.720 -0.400 10.560 0.400 ;
        RECT  9.380 -0.400 9.720 0.575 ;
        RECT  8.190 -0.400 9.380 0.400 ;
        RECT  7.850 -0.400 8.190 0.575 ;
        RECT  5.770 -0.400 7.850 0.400 ;
        RECT  5.430 -0.400 5.770 0.575 ;
        RECT  2.740 -0.400 5.430 0.400 ;
        RECT  2.400 -0.400 2.740 0.575 ;
        RECT  0.520 -0.400 2.400 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.770 4.640 10.560 5.440 ;
        RECT  9.350 4.465 9.770 5.440 ;
        RECT  8.260 4.640 9.350 5.440 ;
        RECT  7.920 4.465 8.260 5.440 ;
        RECT  6.200 4.640 7.920 5.440 ;
        RECT  5.860 4.465 6.200 5.440 ;
        RECT  3.460 4.640 5.860 5.440 ;
        RECT  3.120 4.005 3.460 5.440 ;
        RECT  0.520 4.640 3.120 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.685 2.070 9.740 2.410 ;
        RECT  9.455 0.885 9.685 4.015 ;
        RECT  9.125 0.885 9.455 1.115 ;
        RECT  9.400 2.070 9.455 2.410 ;
        RECT  9.065 3.785 9.455 4.015 ;
        RECT  8.895 0.655 9.125 1.115 ;
        RECT  8.835 3.785 9.065 4.365 ;
        RECT  8.680 0.655 8.895 0.885 ;
        RECT  8.650 4.005 8.835 4.365 ;
        RECT  5.330 4.005 8.650 4.235 ;
        RECT  8.205 2.070 8.540 2.410 ;
        RECT  7.975 2.070 8.205 3.775 ;
        RECT  4.160 3.545 7.975 3.775 ;
        RECT  7.280 0.650 7.510 3.315 ;
        RECT  7.010 0.650 7.280 0.990 ;
        RECT  7.160 2.830 7.280 3.315 ;
        RECT  4.680 3.085 7.160 3.315 ;
        RECT  6.825 1.635 7.035 2.015 ;
        RECT  6.695 1.635 6.825 2.855 ;
        RECT  6.465 0.850 6.695 2.855 ;
        RECT  6.270 0.850 6.465 1.190 ;
        RECT  5.140 2.625 6.465 2.855 ;
        RECT  4.910 1.610 5.140 2.855 ;
        RECT  4.670 1.610 4.910 1.840 ;
        RECT  4.450 2.260 4.680 3.315 ;
        RECT  4.330 1.500 4.670 1.840 ;
        RECT  4.340 2.260 4.450 2.600 ;
        RECT  4.050 0.830 4.390 1.170 ;
        RECT  4.015 1.610 4.330 1.840 ;
        RECT  3.820 3.255 4.160 3.775 ;
        RECT  3.315 0.940 4.050 1.170 ;
        RECT  3.785 1.610 4.015 2.725 ;
        RECT  1.780 3.545 3.820 3.775 ;
        RECT  2.095 2.495 3.785 2.725 ;
        RECT  3.085 0.940 3.315 1.510 ;
        RECT  1.900 1.280 3.085 1.510 ;
        RECT  1.865 2.360 2.095 2.725 ;
        RECT  1.120 0.765 1.930 0.995 ;
        RECT  1.585 1.280 1.900 1.620 ;
        RECT  1.585 3.110 1.780 3.775 ;
        RECT  1.250 4.020 1.590 4.360 ;
        RECT  1.560 1.280 1.585 3.775 ;
        RECT  1.495 1.335 1.560 3.775 ;
        RECT  1.355 1.335 1.495 3.450 ;
        RECT  1.120 4.020 1.250 4.250 ;
        RECT  0.890 0.765 1.120 4.250 ;
        RECT  0.780 1.330 0.890 1.670 ;
        RECT  0.740 3.000 0.890 3.340 ;
    END
END TLATSXL

MACRO TLATSX4
    CLASS CORE ;
    FOREIGN TLATSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.090 0.555 2.430 ;
        RECT  0.140 1.845 0.545 2.430 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.680 1.355 13.060 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.740 1.355 11.760 1.845 ;
        RECT  11.740 2.880 11.760 3.220 ;
        RECT  11.420 1.355 11.740 3.220 ;
        RECT  11.360 1.820 11.420 3.220 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  7.780 1.380 7.865 1.720 ;
        RECT  7.475 1.380 7.780 2.075 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.250 2.070 3.360 2.580 ;
        RECT  3.020 1.845 3.250 2.580 ;
        RECT  2.855 1.845 3.020 2.075 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.680 -0.400 13.860 0.400 ;
        RECT  13.340 -0.400 13.680 0.950 ;
        RECT  12.400 -0.400 13.340 0.400 ;
        RECT  12.060 -0.400 12.400 0.950 ;
        RECT  11.120 -0.400 12.060 0.400 ;
        RECT  10.780 -0.400 11.120 0.950 ;
        RECT  9.700 -0.400 10.780 0.400 ;
        RECT  9.360 -0.400 9.700 1.380 ;
        RECT  7.440 -0.400 9.360 0.400 ;
        RECT  7.100 -0.400 7.440 0.575 ;
        RECT  5.380 -0.400 7.100 0.400 ;
        RECT  5.040 -0.400 5.380 0.575 ;
        RECT  2.700 -0.400 5.040 0.400 ;
        RECT  2.360 -0.400 2.700 0.575 ;
        RECT  0.520 -0.400 2.360 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.680 4.640 13.860 5.440 ;
        RECT  13.340 4.090 13.680 5.440 ;
        RECT  12.400 4.640 13.340 5.440 ;
        RECT  12.060 4.090 12.400 5.440 ;
        RECT  11.080 4.640 12.060 5.440 ;
        RECT  10.740 4.465 11.080 5.440 ;
        RECT  9.840 4.640 10.740 5.440 ;
        RECT  9.500 4.465 9.840 5.440 ;
        RECT  8.020 4.640 9.500 5.440 ;
        RECT  7.680 4.465 8.020 5.440 ;
        RECT  3.620 4.640 7.680 5.440 ;
        RECT  3.280 3.815 3.620 5.440 ;
        RECT  0.520 4.640 3.280 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 2.070 13.670 2.410 ;
        RECT  13.385 2.070 13.615 3.830 ;
        RECT  13.330 2.070 13.385 2.410 ;
        RECT  10.500 3.600 13.385 3.830 ;
        RECT  10.880 1.330 11.110 3.060 ;
        RECT  10.420 1.330 10.880 1.560 ;
        RECT  10.500 2.830 10.880 3.060 ;
        RECT  9.865 2.070 10.650 2.410 ;
        RECT  10.160 2.830 10.500 4.175 ;
        RECT  10.135 1.045 10.420 1.560 ;
        RECT  7.490 3.945 10.160 4.175 ;
        RECT  10.080 1.045 10.135 1.385 ;
        RECT  9.635 2.070 9.865 3.585 ;
        RECT  5.960 3.355 9.635 3.585 ;
        RECT  9.065 2.895 9.180 3.125 ;
        RECT  8.900 1.220 9.065 3.125 ;
        RECT  8.835 1.050 8.900 3.125 ;
        RECT  8.615 1.050 8.835 1.450 ;
        RECT  6.630 2.895 8.835 3.125 ;
        RECT  8.560 1.050 8.615 1.390 ;
        RECT  8.480 1.700 8.535 2.050 ;
        RECT  8.325 1.700 8.480 2.625 ;
        RECT  8.095 0.810 8.325 2.625 ;
        RECT  7.860 0.810 8.095 1.150 ;
        RECT  7.090 2.395 8.095 2.625 ;
        RECT  7.150 3.945 7.490 4.195 ;
        RECT  6.860 1.510 7.090 2.625 ;
        RECT  6.410 1.510 6.860 1.740 ;
        RECT  6.400 2.220 6.630 3.125 ;
        RECT  6.070 1.400 6.410 1.740 ;
        RECT  6.290 2.220 6.400 2.560 ;
        RECT  5.740 0.830 6.080 1.170 ;
        RECT  5.830 1.510 6.070 1.740 ;
        RECT  5.150 3.355 5.960 3.695 ;
        RECT  5.600 1.510 5.830 3.045 ;
        RECT  5.225 0.940 5.740 1.170 ;
        RECT  5.490 2.600 5.600 3.045 ;
        RECT  2.495 2.815 5.490 3.045 ;
        RECT  4.995 0.940 5.225 1.300 ;
        RECT  1.780 3.355 5.150 3.585 ;
        RECT  4.050 1.070 4.995 1.300 ;
        RECT  3.710 0.960 4.050 1.300 ;
        RECT  2.475 1.070 3.710 1.300 ;
        RECT  2.265 2.350 2.495 3.045 ;
        RECT  2.245 1.070 2.475 1.490 ;
        RECT  2.110 2.350 2.265 2.580 ;
        RECT  1.780 1.260 2.245 1.490 ;
        RECT  1.770 2.240 2.110 2.580 ;
        RECT  1.080 0.765 1.930 0.995 ;
        RECT  1.540 1.260 1.780 1.600 ;
        RECT  1.540 3.085 1.780 3.895 ;
        RECT  1.440 1.260 1.540 3.895 ;
        RECT  1.310 1.260 1.440 3.660 ;
        RECT  0.850 0.765 1.080 3.775 ;
        RECT  0.740 1.250 0.850 1.590 ;
        RECT  0.740 2.965 0.850 3.775 ;
    END
END TLATSX4

MACRO TLATSX2
    CLASS CORE ;
    FOREIGN TLATSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.080 0.555 2.420 ;
        RECT  0.140 1.840 0.545 2.420 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.005 2.630 11.040 4.255 ;
        RECT  11.005 0.765 11.025 1.575 ;
        RECT  10.775 0.765 11.005 4.255 ;
        RECT  10.685 0.765 10.775 1.575 ;
        RECT  10.700 2.630 10.775 4.255 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.765 1.445 9.995 3.050 ;
        RECT  9.400 1.445 9.765 1.675 ;
        RECT  9.600 2.820 9.765 3.050 ;
        RECT  9.260 2.820 9.600 3.195 ;
        RECT  9.060 1.335 9.400 1.675 ;
        RECT  8.795 2.935 9.260 3.195 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 1.500 6.130 1.840 ;
        RECT  5.725 1.500 5.790 1.730 ;
        RECT  5.495 1.285 5.725 1.730 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 1.795 3.395 2.200 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.220 -0.400 11.220 0.400 ;
        RECT  9.880 -0.400 10.220 0.575 ;
        RECT  7.960 -0.400 9.880 0.400 ;
        RECT  7.620 -0.400 7.960 1.210 ;
        RECT  5.660 -0.400 7.620 0.400 ;
        RECT  5.320 -0.400 5.660 0.575 ;
        RECT  2.880 -0.400 5.320 0.400 ;
        RECT  2.540 -0.400 2.880 0.575 ;
        RECT  0.520 -0.400 2.540 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 4.640 11.220 5.440 ;
        RECT  9.980 4.080 10.320 5.440 ;
        RECT  8.200 4.640 9.980 5.440 ;
        RECT  7.860 4.465 8.200 5.440 ;
        RECT  6.200 4.640 7.860 5.440 ;
        RECT  5.860 4.465 6.200 5.440 ;
        RECT  3.700 4.640 5.860 5.440 ;
        RECT  3.360 4.090 3.700 5.440 ;
        RECT  0.520 4.640 3.360 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.225 0.870 10.455 3.850 ;
        RECT  8.680 0.870 10.225 1.100 ;
        RECT  8.985 3.620 10.225 3.850 ;
        RECT  8.205 2.070 9.060 2.410 ;
        RECT  8.620 3.620 8.985 4.175 ;
        RECT  8.340 0.870 8.680 1.210 ;
        RECT  5.670 3.945 8.620 4.175 ;
        RECT  7.975 2.070 8.205 3.655 ;
        RECT  1.820 3.425 7.975 3.655 ;
        RECT  7.390 2.855 7.500 3.195 ;
        RECT  7.160 0.980 7.390 3.195 ;
        RECT  6.820 0.870 7.160 1.210 ;
        RECT  4.650 2.965 7.160 3.195 ;
        RECT  6.825 1.605 6.915 1.975 ;
        RECT  6.590 1.605 6.825 2.735 ;
        RECT  6.360 0.850 6.590 2.735 ;
        RECT  6.120 0.850 6.360 1.190 ;
        RECT  5.110 2.505 6.360 2.735 ;
        RECT  5.330 3.945 5.670 4.225 ;
        RECT  4.880 1.890 5.110 2.735 ;
        RECT  4.650 1.890 4.880 2.120 ;
        RECT  4.310 1.780 4.650 2.120 ;
        RECT  4.420 2.505 4.650 3.195 ;
        RECT  4.230 2.505 4.420 2.735 ;
        RECT  3.925 1.890 4.310 2.120 ;
        RECT  4.190 0.810 4.300 1.150 ;
        RECT  3.960 0.810 4.190 1.490 ;
        RECT  1.900 1.260 3.960 1.490 ;
        RECT  3.695 1.890 3.925 3.195 ;
        RECT  2.475 2.965 3.695 3.195 ;
        RECT  2.245 2.230 2.475 3.195 ;
        RECT  2.190 2.230 2.245 2.460 ;
        RECT  1.850 2.120 2.190 2.460 ;
        RECT  1.120 0.765 1.930 0.995 ;
        RECT  1.620 1.260 1.900 1.600 ;
        RECT  1.620 3.080 1.820 3.890 ;
        RECT  1.480 1.260 1.620 3.890 ;
        RECT  1.390 1.260 1.480 3.655 ;
        RECT  0.890 0.765 1.120 3.120 ;
        RECT  0.780 1.290 0.890 1.630 ;
        RECT  0.780 2.780 0.890 3.120 ;
    END
END TLATSX2

MACRO TLATSX1
    CLASS CORE ;
    FOREIGN TLATSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 2.015 0.560 2.355 ;
        RECT  0.140 1.820 0.550 2.355 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 1.320 10.360 1.845 ;
        RECT  10.345 3.020 10.360 3.360 ;
        RECT  10.115 1.320 10.345 3.360 ;
        RECT  10.040 1.320 10.115 1.845 ;
        RECT  10.020 3.020 10.115 3.360 ;
        RECT  10.020 1.320 10.040 1.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.925 1.430 9.155 3.310 ;
        RECT  8.640 1.430 8.925 1.770 ;
        RECT  8.680 2.940 8.925 3.310 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.890 1.500 6.230 1.840 ;
        RECT  5.725 1.500 5.890 1.730 ;
        RECT  5.495 1.285 5.725 1.730 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.830 1.845 3.460 2.185 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.720 -0.400 10.560 0.400 ;
        RECT  9.380 -0.400 9.720 0.575 ;
        RECT  8.170 -0.400 9.380 0.400 ;
        RECT  7.830 -0.400 8.170 0.575 ;
        RECT  5.770 -0.400 7.830 0.400 ;
        RECT  5.430 -0.400 5.770 0.575 ;
        RECT  2.740 -0.400 5.430 0.400 ;
        RECT  2.400 -0.400 2.740 0.575 ;
        RECT  0.520 -0.400 2.400 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.775 4.640 10.560 5.440 ;
        RECT  9.350 4.465 9.775 5.440 ;
        RECT  8.260 4.640 9.350 5.440 ;
        RECT  7.920 4.465 8.260 5.440 ;
        RECT  6.200 4.640 7.920 5.440 ;
        RECT  5.860 4.465 6.200 5.440 ;
        RECT  3.460 4.640 5.860 5.440 ;
        RECT  3.120 4.080 3.460 5.440 ;
        RECT  0.520 4.640 3.120 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.455 0.885 9.685 4.015 ;
        RECT  9.125 0.885 9.455 1.115 ;
        RECT  9.040 3.785 9.455 4.015 ;
        RECT  8.895 0.675 9.125 1.115 ;
        RECT  8.810 3.785 9.040 4.365 ;
        RECT  8.680 0.675 8.895 0.905 ;
        RECT  8.680 4.005 8.810 4.365 ;
        RECT  5.330 4.005 8.680 4.235 ;
        RECT  8.205 2.070 8.540 2.410 ;
        RECT  7.975 2.070 8.205 3.775 ;
        RECT  4.160 3.545 7.975 3.775 ;
        RECT  7.445 1.020 7.500 3.170 ;
        RECT  7.270 1.020 7.445 3.315 ;
        RECT  7.010 1.020 7.270 1.360 ;
        RECT  7.160 2.830 7.270 3.315 ;
        RECT  4.680 3.085 7.160 3.315 ;
        RECT  6.825 1.635 7.035 2.015 ;
        RECT  6.695 1.635 6.825 2.855 ;
        RECT  6.465 0.850 6.695 2.855 ;
        RECT  6.270 0.850 6.465 1.190 ;
        RECT  5.140 2.625 6.465 2.855 ;
        RECT  4.910 1.610 5.140 2.855 ;
        RECT  4.670 1.610 4.910 1.840 ;
        RECT  4.450 2.260 4.680 3.315 ;
        RECT  4.330 1.500 4.670 1.840 ;
        RECT  4.340 2.260 4.450 2.600 ;
        RECT  4.030 0.810 4.370 1.150 ;
        RECT  4.015 1.610 4.330 1.840 ;
        RECT  3.820 3.490 4.160 3.830 ;
        RECT  3.315 0.920 4.030 1.150 ;
        RECT  3.785 1.610 4.015 2.725 ;
        RECT  1.780 3.545 3.820 3.775 ;
        RECT  2.095 2.495 3.785 2.725 ;
        RECT  3.085 0.920 3.315 1.565 ;
        RECT  1.585 1.335 3.085 1.565 ;
        RECT  1.865 2.360 2.095 2.725 ;
        RECT  1.120 0.765 1.930 0.995 ;
        RECT  1.585 3.110 1.780 3.775 ;
        RECT  1.250 4.020 1.590 4.360 ;
        RECT  1.495 1.335 1.585 3.775 ;
        RECT  1.355 1.335 1.495 3.450 ;
        RECT  1.120 4.020 1.250 4.250 ;
        RECT  0.890 0.765 1.120 4.250 ;
        RECT  0.780 1.330 0.890 1.670 ;
        RECT  0.740 2.980 0.890 3.320 ;
    END
END TLATSX1

MACRO TLATRXL
    CLASS CORE ;
    FOREIGN TLATRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.710 2.090 4.850 2.320 ;
        RECT  4.480 2.090 4.710 2.885 ;
        RECT  4.175 2.405 4.480 2.885 ;
        RECT  3.745 2.655 4.175 2.885 ;
        RECT  3.405 2.655 3.745 3.130 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.365 1.230 8.400 1.570 ;
        RECT  8.365 3.050 8.400 3.390 ;
        RECT  8.135 1.230 8.365 3.390 ;
        RECT  8.060 1.230 8.135 1.570 ;
        RECT  8.060 3.050 8.135 3.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.505 0.810 7.735 3.755 ;
        RECT  6.960 0.810 7.505 1.040 ;
        RECT  7.140 3.525 7.505 3.755 ;
        RECT  6.800 3.525 7.140 4.140 ;
        RECT  6.620 0.700 6.960 1.040 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.840 0.530 2.490 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.405 2.425 3.075 ;
        RECT  1.995 2.735 2.120 3.075 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.720 -0.400 8.580 0.400 ;
        RECT  7.380 -0.400 7.720 0.575 ;
        RECT  6.080 -0.400 7.380 0.400 ;
        RECT  5.740 -0.400 6.080 0.575 ;
        RECT  2.020 -0.400 5.740 0.400 ;
        RECT  1.680 -0.400 2.020 0.575 ;
        RECT  0.520 -0.400 1.680 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.840 4.640 8.580 5.440 ;
        RECT  7.500 4.465 7.840 5.440 ;
        RECT  6.380 4.640 7.500 5.440 ;
        RECT  6.040 4.465 6.380 5.440 ;
        RECT  4.175 4.640 6.040 5.440 ;
        RECT  3.835 3.850 4.175 5.440 ;
        RECT  2.095 4.640 3.835 5.440 ;
        RECT  1.755 3.570 2.095 5.440 ;
        RECT  0.520 4.640 1.755 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.045 1.600 7.275 3.175 ;
        RECT  6.960 1.600 7.045 1.830 ;
        RECT  6.800 2.810 7.045 3.175 ;
        RECT  6.620 1.490 6.960 1.830 ;
        RECT  6.395 2.945 6.800 3.175 ;
        RECT  6.320 2.070 6.660 2.410 ;
        RECT  6.165 2.945 6.395 4.195 ;
        RECT  5.835 2.125 6.320 2.355 ;
        RECT  5.480 3.965 6.165 4.195 ;
        RECT  5.825 2.125 5.835 3.510 ;
        RECT  5.605 1.170 5.825 3.510 ;
        RECT  5.595 1.170 5.605 2.355 ;
        RECT  4.935 3.280 5.605 3.510 ;
        RECT  3.900 1.170 5.595 1.400 ;
        RECT  5.080 1.630 5.310 3.045 ;
        RECT  3.660 1.630 5.080 1.860 ;
        RECT  4.940 2.705 5.080 3.045 ;
        RECT  4.570 3.280 4.935 3.620 ;
        RECT  3.375 3.390 4.570 3.620 ;
        RECT  3.560 1.060 3.900 1.400 ;
        RECT  3.320 1.630 3.660 1.970 ;
        RECT  3.035 3.390 3.375 3.770 ;
        RECT  1.675 1.685 3.320 1.915 ;
        RECT  1.525 0.810 1.675 3.175 ;
        RECT  1.445 0.810 1.525 3.910 ;
        RECT  1.220 0.810 1.445 1.040 ;
        RECT  1.295 2.945 1.445 3.910 ;
        RECT  1.035 3.570 1.295 3.910 ;
        RECT  0.880 0.700 1.220 1.040 ;
        RECT  1.065 2.270 1.215 2.610 ;
        RECT  1.065 1.400 1.120 1.740 ;
        RECT  0.835 1.400 1.065 3.190 ;
        RECT  0.780 1.400 0.835 1.740 ;
    END
END TLATRXL

MACRO TLATRX4
    CLASS CORE ;
    FOREIGN TLATRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 2.720 3.270 3.060 ;
        RECT  2.855 2.405 3.160 3.060 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.060 1.820 11.080 3.220 ;
        RECT  10.720 1.455 11.060 3.220 ;
        RECT  10.700 1.820 10.720 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.760 1.455 9.780 1.845 ;
        RECT  9.760 2.635 9.780 3.180 ;
        RECT  9.440 1.455 9.760 3.220 ;
        RECT  9.380 1.820 9.440 3.220 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 2.045 6.350 2.275 ;
        RECT  6.065 1.845 6.295 2.275 ;
        RECT  5.715 1.845 6.065 2.270 ;
        RECT  5.495 1.845 5.715 2.075 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 1.820 2.090 2.340 ;
        RECT  1.460 1.820 1.750 2.180 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.700 -0.400 11.880 0.400 ;
        RECT  11.360 -0.400 11.700 1.045 ;
        RECT  10.420 -0.400 11.360 0.400 ;
        RECT  10.080 -0.400 10.420 1.045 ;
        RECT  9.060 -0.400 10.080 0.400 ;
        RECT  8.720 -0.400 9.060 0.575 ;
        RECT  7.800 -0.400 8.720 0.400 ;
        RECT  7.460 -0.400 7.800 0.575 ;
        RECT  6.200 -0.400 7.460 0.400 ;
        RECT  5.860 -0.400 6.200 0.575 ;
        RECT  2.440 -0.400 5.860 0.400 ;
        RECT  2.100 -0.400 2.440 1.055 ;
        RECT  0.000 -0.400 2.100 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.700 4.640 11.880 5.440 ;
        RECT  11.360 4.090 11.700 5.440 ;
        RECT  10.420 4.640 11.360 5.440 ;
        RECT  10.080 4.090 10.420 5.440 ;
        RECT  9.095 4.640 10.080 5.440 ;
        RECT  8.675 4.465 9.095 5.440 ;
        RECT  7.620 4.640 8.675 5.440 ;
        RECT  7.280 4.465 7.620 5.440 ;
        RECT  5.360 4.640 7.280 5.440 ;
        RECT  5.020 4.465 5.360 5.440 ;
        RECT  3.120 4.640 5.020 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  0.520 4.640 2.780 5.440 ;
        RECT  0.180 4.145 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.385 2.100 11.615 3.860 ;
        RECT  8.865 3.630 11.385 3.860 ;
        RECT  8.635 1.565 8.865 3.860 ;
        RECT  8.500 1.565 8.635 1.795 ;
        RECT  8.375 3.630 8.635 3.860 ;
        RECT  8.160 1.455 8.500 1.795 ;
        RECT  8.145 3.035 8.375 4.175 ;
        RECT  8.000 2.200 8.340 2.540 ;
        RECT  4.775 3.945 8.145 4.175 ;
        RECT  7.915 2.310 8.000 2.540 ;
        RECT  7.685 2.310 7.915 3.655 ;
        RECT  7.455 1.090 7.800 1.430 ;
        RECT  3.920 3.425 7.685 3.655 ;
        RECT  7.225 0.805 7.455 3.195 ;
        RECT  5.165 0.805 7.225 1.035 ;
        RECT  6.520 2.965 7.225 3.195 ;
        RECT  6.765 1.410 6.995 2.735 ;
        RECT  6.570 1.410 6.765 1.750 ;
        RECT  6.160 2.505 6.765 2.735 ;
        RECT  5.930 2.505 6.160 3.135 ;
        RECT  4.675 2.905 5.930 3.135 ;
        RECT  4.935 0.805 5.165 2.450 ;
        RECT  4.300 2.220 4.935 2.450 ;
        RECT  4.545 3.945 4.775 4.310 ;
        RECT  4.350 1.550 4.690 1.975 ;
        RECT  4.445 2.790 4.675 3.135 ;
        RECT  3.730 2.790 4.445 3.020 ;
        RECT  3.730 1.745 4.350 1.975 ;
        RECT  4.115 0.980 4.320 1.320 ;
        RECT  3.960 2.220 4.300 2.560 ;
        RECT  3.820 3.970 4.160 4.310 ;
        RECT  3.885 0.980 4.115 1.515 ;
        RECT  3.580 3.290 3.920 3.655 ;
        RECT  1.035 1.285 3.885 1.515 ;
        RECT  1.125 3.970 3.820 4.200 ;
        RECT  3.500 1.745 3.730 3.020 ;
        RECT  1.800 3.425 3.580 3.655 ;
        RECT  2.550 1.745 3.500 1.975 ;
        RECT  2.320 1.745 2.550 2.970 ;
        RECT  1.460 2.740 2.320 2.970 ;
        RECT  1.690 3.315 1.800 3.655 ;
        RECT  1.460 3.220 1.690 3.655 ;
        RECT  1.035 3.220 1.460 3.450 ;
        RECT  0.895 3.685 1.125 4.200 ;
        RECT  0.805 1.285 1.035 3.450 ;
        RECT  0.495 3.685 0.895 3.915 ;
        RECT  0.520 1.285 0.805 1.515 ;
        RECT  0.495 1.835 0.550 2.175 ;
        RECT  0.180 1.120 0.520 1.515 ;
        RECT  0.265 1.835 0.495 3.915 ;
        RECT  0.210 1.835 0.265 2.175 ;
    END
END TLATRX4

MACRO TLATRX2
    CLASS CORE ;
    FOREIGN TLATRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATRXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.135 2.940 4.475 3.510 ;
        RECT  3.390 2.940 4.135 3.170 ;
        RECT  3.160 2.310 3.390 3.170 ;
        RECT  3.030 2.310 3.160 2.540 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.720 0.775 9.060 4.275 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.540 2.965 7.705 3.195 ;
        RECT  7.200 1.390 7.540 4.110 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.845 0.530 2.525 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.275 2.700 2.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 -0.400 9.240 0.400 ;
        RECT  7.960 -0.400 8.300 0.575 ;
        RECT  6.080 -0.400 7.960 0.400 ;
        RECT  5.740 -0.400 6.080 0.575 ;
        RECT  2.420 -0.400 5.740 0.400 ;
        RECT  2.080 -0.400 2.420 0.575 ;
        RECT  0.520 -0.400 2.080 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 4.640 9.240 5.440 ;
        RECT  7.960 3.910 8.300 5.440 ;
        RECT  6.270 4.640 7.960 5.440 ;
        RECT  5.855 4.465 6.270 5.440 ;
        RECT  4.200 4.640 5.855 5.440 ;
        RECT  3.860 4.465 4.200 5.440 ;
        RECT  2.120 4.640 3.860 5.440 ;
        RECT  1.780 4.090 2.120 5.440 ;
        RECT  0.520 4.640 1.780 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.340 2.100 8.450 2.440 ;
        RECT  8.110 0.865 8.340 2.440 ;
        RECT  6.840 0.865 8.110 1.095 ;
        RECT  6.785 0.865 6.840 1.410 ;
        RECT  6.785 3.440 6.840 3.780 ;
        RECT  6.555 0.865 6.785 3.780 ;
        RECT  6.500 0.865 6.555 1.410 ;
        RECT  6.060 2.030 6.555 2.370 ;
        RECT  6.500 3.440 6.555 3.780 ;
        RECT  5.725 2.705 6.315 3.050 ;
        RECT  5.495 0.890 5.725 4.135 ;
        RECT  4.300 0.890 5.495 1.120 ;
        RECT  3.400 3.905 5.495 4.135 ;
        RECT  5.070 3.295 5.180 3.635 ;
        RECT  4.840 2.330 5.070 3.635 ;
        RECT  4.040 2.330 4.840 2.560 ;
        RECT  4.600 1.760 4.710 2.100 ;
        RECT  4.370 1.350 4.600 2.100 ;
        RECT  2.525 1.350 4.370 1.580 ;
        RECT  3.960 0.780 4.300 1.120 ;
        RECT  3.810 1.815 4.040 2.560 ;
        RECT  1.825 1.815 3.810 2.045 ;
        RECT  3.060 3.770 3.400 4.135 ;
        RECT  2.295 0.820 2.525 1.580 ;
        RECT  1.120 0.820 2.295 1.050 ;
        RECT  1.675 1.295 1.825 2.045 ;
        RECT  1.445 1.295 1.675 3.860 ;
        RECT  1.300 3.630 1.445 3.860 ;
        RECT  0.960 3.630 1.300 3.970 ;
        RECT  1.120 2.060 1.215 2.405 ;
        RECT  0.890 0.820 1.120 3.120 ;
        RECT  0.780 1.240 0.890 1.580 ;
        RECT  0.780 2.780 0.890 3.120 ;
    END
END TLATRX2

MACRO TLATRX1
    CLASS CORE ;
    FOREIGN TLATRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATRXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.710 2.000 4.850 2.230 ;
        RECT  4.480 2.000 4.710 2.635 ;
        RECT  3.745 2.405 4.480 2.635 ;
        RECT  3.515 2.405 3.745 3.130 ;
        RECT  3.405 2.630 3.515 3.130 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 1.200 8.400 3.300 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.505 0.865 7.735 3.755 ;
        RECT  6.960 0.865 7.505 1.095 ;
        RECT  7.075 3.525 7.505 3.755 ;
        RECT  6.845 3.525 7.075 4.010 ;
        RECT  6.620 0.700 6.960 1.095 ;
        RECT  6.815 3.525 6.845 3.755 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.845 0.530 2.475 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.405 2.425 3.095 ;
        RECT  1.995 2.755 2.120 3.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.720 -0.400 8.580 0.400 ;
        RECT  7.380 -0.400 7.720 0.575 ;
        RECT  6.080 -0.400 7.380 0.400 ;
        RECT  5.740 -0.400 6.080 0.575 ;
        RECT  2.020 -0.400 5.740 0.400 ;
        RECT  1.680 -0.400 2.020 0.575 ;
        RECT  0.520 -0.400 1.680 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.730 4.640 8.580 5.440 ;
        RECT  7.305 4.465 7.730 5.440 ;
        RECT  6.370 4.640 7.305 5.440 ;
        RECT  6.030 4.465 6.370 5.440 ;
        RECT  4.175 4.640 6.030 5.440 ;
        RECT  3.835 3.850 4.175 5.440 ;
        RECT  2.095 4.640 3.835 5.440 ;
        RECT  1.755 3.620 2.095 5.440 ;
        RECT  0.520 4.640 1.755 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.045 1.600 7.275 3.175 ;
        RECT  6.960 1.600 7.045 1.830 ;
        RECT  6.790 2.810 7.045 3.175 ;
        RECT  6.620 1.490 6.960 1.830 ;
        RECT  6.395 2.945 6.790 3.175 ;
        RECT  6.320 2.070 6.660 2.410 ;
        RECT  6.165 2.945 6.395 4.125 ;
        RECT  5.835 2.125 6.320 2.355 ;
        RECT  5.480 3.895 6.165 4.125 ;
        RECT  5.825 2.125 5.835 3.460 ;
        RECT  5.605 1.070 5.825 3.460 ;
        RECT  5.595 1.070 5.605 2.355 ;
        RECT  4.935 3.230 5.605 3.460 ;
        RECT  3.900 1.070 5.595 1.300 ;
        RECT  5.080 1.530 5.310 2.955 ;
        RECT  3.660 1.530 5.080 1.760 ;
        RECT  4.940 2.615 5.080 2.955 ;
        RECT  4.570 3.230 4.935 3.620 ;
        RECT  3.375 3.390 4.570 3.620 ;
        RECT  3.560 0.960 3.900 1.300 ;
        RECT  3.320 1.530 3.660 1.950 ;
        RECT  3.035 3.390 3.375 3.730 ;
        RECT  1.675 1.665 3.320 1.895 ;
        RECT  1.525 0.810 1.675 3.175 ;
        RECT  1.445 0.810 1.525 3.960 ;
        RECT  1.220 0.810 1.445 1.040 ;
        RECT  1.295 2.945 1.445 3.960 ;
        RECT  1.035 3.620 1.295 3.960 ;
        RECT  0.880 0.700 1.220 1.040 ;
        RECT  1.065 2.270 1.215 2.610 ;
        RECT  0.835 1.400 1.065 3.190 ;
    END
END TLATRX1

MACRO TLATNSRXL
    CLASS CORE ;
    FOREIGN TLATNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.105 0.555 2.445 ;
        RECT  0.140 1.840 0.545 2.445 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.510 1.820 3.845 2.600 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.005 1.240 11.040 1.580 ;
        RECT  11.005 3.020 11.040 3.360 ;
        RECT  10.775 1.240 11.005 3.360 ;
        RECT  10.700 1.240 10.775 1.580 ;
        RECT  10.700 3.020 10.775 3.360 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.640 2.965 9.685 3.205 ;
        RECT  9.620 2.965 9.640 3.310 ;
        RECT  9.390 1.430 9.620 3.310 ;
        RECT  9.280 1.430 9.390 1.770 ;
        RECT  9.300 2.970 9.390 3.310 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 1.930 6.900 2.270 ;
        RECT  6.385 1.930 6.560 2.160 ;
        RECT  6.155 1.845 6.385 2.160 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.900 3.085 2.660 ;
        RECT  2.580 1.900 2.780 2.240 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 -0.400 11.220 0.400 ;
        RECT  9.980 -0.400 10.320 0.575 ;
        RECT  8.820 -0.400 9.980 0.400 ;
        RECT  8.480 -0.400 8.820 0.575 ;
        RECT  6.690 -0.400 8.480 0.400 ;
        RECT  6.350 -0.400 6.690 0.575 ;
        RECT  2.720 -0.400 6.350 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  0.520 -0.400 2.380 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 4.640 11.220 5.440 ;
        RECT  9.970 4.465 10.405 5.440 ;
        RECT  8.880 4.640 9.970 5.440 ;
        RECT  8.540 4.465 8.880 5.440 ;
        RECT  6.820 4.640 8.540 5.440 ;
        RECT  6.480 4.465 6.820 5.440 ;
        RECT  3.500 4.640 6.480 5.440 ;
        RECT  3.160 4.135 3.500 5.440 ;
        RECT  0.520 4.640 3.160 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.415 2.070 10.470 2.410 ;
        RECT  10.185 0.805 10.415 4.015 ;
        RECT  9.620 0.805 10.185 1.035 ;
        RECT  10.130 2.070 10.185 2.410 ;
        RECT  9.640 3.785 10.185 4.015 ;
        RECT  9.410 3.785 9.640 4.365 ;
        RECT  9.280 0.635 9.620 1.035 ;
        RECT  9.300 4.005 9.410 4.365 ;
        RECT  5.950 4.005 9.300 4.235 ;
        RECT  9.025 2.090 9.160 2.430 ;
        RECT  8.795 2.090 9.025 3.775 ;
        RECT  4.765 3.545 8.795 3.775 ;
        RECT  7.965 0.745 8.195 3.270 ;
        RECT  7.680 0.745 7.965 1.085 ;
        RECT  7.780 2.930 7.965 3.270 ;
        RECT  7.485 1.900 7.730 2.240 ;
        RECT  5.655 0.855 7.680 1.085 ;
        RECT  7.255 1.315 7.485 3.315 ;
        RECT  6.980 1.315 7.255 1.545 ;
        RECT  5.585 3.085 7.255 3.315 ;
        RECT  5.425 0.855 5.655 1.940 ;
        RECT  5.355 2.490 5.585 3.315 ;
        RECT  5.010 1.710 5.425 1.940 ;
        RECT  5.190 2.490 5.355 2.720 ;
        RECT  4.850 2.380 5.190 2.720 ;
        RECT  4.670 1.710 5.010 2.050 ;
        RECT  4.535 3.210 4.765 3.775 ;
        RECT  4.305 1.820 4.670 2.050 ;
        RECT  4.260 1.130 4.600 1.470 ;
        RECT  1.820 3.545 4.535 3.775 ;
        RECT  4.075 1.820 4.305 3.120 ;
        RECT  2.595 1.240 4.260 1.470 ;
        RECT  2.475 2.890 4.075 3.120 ;
        RECT  2.365 1.240 2.595 1.545 ;
        RECT  2.245 2.470 2.475 3.120 ;
        RECT  1.620 1.315 2.365 1.545 ;
        RECT  2.190 2.470 2.245 2.700 ;
        RECT  1.850 2.360 2.190 2.700 ;
        RECT  1.620 0.730 1.960 1.070 ;
        RECT  1.620 3.110 1.820 3.775 ;
        RECT  1.290 4.020 1.630 4.360 ;
        RECT  1.120 0.840 1.620 1.070 ;
        RECT  1.590 1.315 1.620 3.775 ;
        RECT  1.390 1.315 1.590 3.450 ;
        RECT  1.120 4.020 1.290 4.250 ;
        RECT  0.890 0.840 1.120 4.250 ;
        RECT  0.780 1.290 0.890 1.630 ;
        RECT  0.780 3.000 0.890 3.340 ;
    END
END TLATNSRXL

MACRO TLATNSRX4
    CLASS CORE ;
    FOREIGN TLATNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.790 1.900 1.105 2.635 ;
        RECT  0.710 1.900 0.790 2.405 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.760 1.735 9.100 2.355 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.680 1.820 15.700 3.220 ;
        RECT  15.340 1.260 15.680 3.220 ;
        RECT  15.320 1.820 15.340 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.380 1.260 14.400 1.600 ;
        RECT  14.380 2.880 14.400 3.220 ;
        RECT  14.060 1.260 14.380 3.220 ;
        RECT  14.000 1.820 14.060 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  10.080 1.490 10.420 2.100 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.950 2.295 5.290 2.635 ;
        RECT  3.745 2.350 4.950 2.580 ;
        RECT  3.515 1.845 3.745 2.580 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 -0.400 16.500 0.400 ;
        RECT  15.980 -0.400 16.320 0.950 ;
        RECT  15.040 -0.400 15.980 0.400 ;
        RECT  14.700 -0.400 15.040 0.950 ;
        RECT  13.720 -0.400 14.700 0.400 ;
        RECT  13.380 -0.400 13.720 0.575 ;
        RECT  12.060 -0.400 13.380 0.400 ;
        RECT  11.720 -0.400 12.060 0.575 ;
        RECT  9.940 -0.400 11.720 0.400 ;
        RECT  9.600 -0.400 9.940 0.575 ;
        RECT  6.100 -0.400 9.600 0.400 ;
        RECT  5.760 -0.400 6.100 0.920 ;
        RECT  2.965 -0.400 5.760 0.400 ;
        RECT  2.625 -0.400 2.965 0.575 ;
        RECT  1.280 -0.400 2.625 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 4.640 16.500 5.440 ;
        RECT  15.980 4.090 16.320 5.440 ;
        RECT  15.040 4.640 15.980 5.440 ;
        RECT  14.700 4.090 15.040 5.440 ;
        RECT  13.720 4.640 14.700 5.440 ;
        RECT  13.380 4.465 13.720 5.440 ;
        RECT  12.160 4.640 13.380 5.440 ;
        RECT  11.820 4.465 12.160 5.440 ;
        RECT  10.340 4.640 11.820 5.440 ;
        RECT  10.000 4.465 10.340 5.440 ;
        RECT  6.980 4.640 10.000 5.440 ;
        RECT  6.640 4.465 6.980 5.440 ;
        RECT  1.240 4.640 6.640 5.440 ;
        RECT  0.900 3.740 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.160 2.070 16.270 2.410 ;
        RECT  15.930 2.070 16.160 3.785 ;
        RECT  12.905 3.555 15.930 3.785 ;
        RECT  13.465 1.370 13.695 3.015 ;
        RECT  12.970 1.370 13.465 1.600 ;
        RECT  12.905 2.785 13.465 3.015 ;
        RECT  12.395 2.080 13.190 2.420 ;
        RECT  12.630 1.260 12.970 1.600 ;
        RECT  12.675 2.785 12.905 4.225 ;
        RECT  9.470 3.995 12.675 4.225 ;
        RECT  12.165 2.080 12.395 3.655 ;
        RECT  2.545 3.425 12.165 3.655 ;
        RECT  11.645 1.225 11.875 3.195 ;
        RECT  11.450 1.225 11.645 1.455 ;
        RECT  8.375 2.965 11.645 3.195 ;
        RECT  11.110 1.115 11.450 1.455 ;
        RECT  10.880 1.685 11.355 2.075 ;
        RECT  10.880 2.505 10.955 2.735 ;
        RECT  10.650 0.810 10.880 2.735 ;
        RECT  10.360 0.810 10.650 1.150 ;
        RECT  10.600 2.505 10.650 2.735 ;
        RECT  8.595 0.865 10.360 1.095 ;
        RECT  7.685 4.180 9.140 4.410 ;
        RECT  8.365 0.865 8.595 1.355 ;
        RECT  8.375 1.585 8.430 1.925 ;
        RECT  8.145 1.585 8.375 3.195 ;
        RECT  7.745 1.125 8.365 1.355 ;
        RECT  8.090 1.585 8.145 1.925 ;
        RECT  3.130 2.965 8.145 3.195 ;
        RECT  6.985 0.665 8.020 0.895 ;
        RECT  7.720 1.125 7.745 2.300 ;
        RECT  7.515 1.125 7.720 2.355 ;
        RECT  7.455 3.945 7.685 4.410 ;
        RECT  7.380 1.835 7.515 2.355 ;
        RECT  6.065 3.945 7.455 4.175 ;
        RECT  7.355 1.835 7.380 2.300 ;
        RECT  4.550 1.835 7.355 2.065 ;
        RECT  6.755 0.665 6.985 1.385 ;
        RECT  4.070 1.155 6.755 1.385 ;
        RECT  5.835 3.945 6.065 4.355 ;
        RECT  1.865 4.125 5.835 4.355 ;
        RECT  4.210 1.780 4.550 2.120 ;
        RECT  3.730 1.100 4.070 1.440 ;
        RECT  2.545 1.155 3.730 1.385 ;
        RECT  2.900 2.210 3.130 3.195 ;
        RECT  2.790 2.210 2.900 2.550 ;
        RECT  2.315 1.155 2.545 3.655 ;
        RECT  1.800 1.155 2.315 1.495 ;
        RECT  1.865 1.790 2.000 2.130 ;
        RECT  1.635 1.790 1.865 4.355 ;
        RECT  1.565 1.790 1.635 2.020 ;
        RECT  0.520 2.980 1.635 3.210 ;
        RECT  1.335 1.180 1.565 2.020 ;
        RECT  0.520 1.180 1.335 1.410 ;
        RECT  0.180 1.070 0.520 1.410 ;
        RECT  0.180 2.980 0.520 3.920 ;
    END
END TLATNSRX4

MACRO TLATNSRX2
    CLASS CORE ;
    FOREIGN TLATNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 2.170 0.560 2.510 ;
        RECT  0.215 1.845 0.550 2.510 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 1.845 4.405 2.100 ;
        RECT  3.650 1.845 3.990 2.330 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 0.765 11.700 1.575 ;
        RECT  11.665 2.975 11.700 4.255 ;
        RECT  11.435 0.765 11.665 4.255 ;
        RECT  11.360 0.765 11.435 1.575 ;
        RECT  11.360 2.975 11.435 4.255 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.260 2.965 10.345 3.195 ;
        RECT  10.180 2.635 10.260 3.195 ;
        RECT  9.975 1.360 10.180 3.195 ;
        RECT  9.950 1.360 9.975 3.180 ;
        RECT  9.840 1.360 9.950 1.700 ;
        RECT  9.920 2.840 9.950 3.180 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.655 2.320 6.930 2.660 ;
        RECT  6.425 1.845 6.655 2.660 ;
        RECT  6.155 1.845 6.425 2.075 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.980 1.845 3.320 2.445 ;
        RECT  2.855 1.845 2.980 2.075 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.940 -0.400 11.880 0.400 ;
        RECT  10.600 -0.400 10.940 0.575 ;
        RECT  8.820 -0.400 10.600 0.400 ;
        RECT  8.480 -0.400 8.820 0.575 ;
        RECT  6.780 -0.400 8.480 0.400 ;
        RECT  6.440 -0.400 6.780 0.575 ;
        RECT  2.830 -0.400 6.440 0.400 ;
        RECT  2.490 -0.400 2.830 0.575 ;
        RECT  0.520 -0.400 2.490 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.980 4.640 11.880 5.440 ;
        RECT  10.640 4.090 10.980 5.440 ;
        RECT  8.800 4.640 10.640 5.440 ;
        RECT  8.460 4.465 8.800 5.440 ;
        RECT  6.900 4.640 8.460 5.440 ;
        RECT  6.560 4.465 6.900 5.440 ;
        RECT  3.620 4.640 6.560 5.440 ;
        RECT  3.280 3.740 3.620 5.440 ;
        RECT  0.520 4.640 3.280 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.900 0.885 11.130 3.835 ;
        RECT  9.480 0.885 10.900 1.115 ;
        RECT  9.560 3.605 10.900 3.835 ;
        RECT  9.220 2.070 9.560 2.410 ;
        RECT  9.450 2.945 9.560 3.835 ;
        RECT  9.140 0.885 9.480 1.430 ;
        RECT  9.220 2.945 9.450 4.235 ;
        RECT  8.765 2.180 9.220 2.410 ;
        RECT  6.030 4.005 9.220 4.235 ;
        RECT  8.535 2.180 8.765 3.655 ;
        RECT  4.900 3.425 8.535 3.655 ;
        RECT  8.065 1.095 8.245 3.190 ;
        RECT  8.015 0.875 8.065 3.190 ;
        RECT  7.780 0.875 8.015 1.440 ;
        RECT  7.860 2.850 8.015 3.190 ;
        RECT  5.755 0.875 7.780 1.105 ;
        RECT  7.500 1.930 7.780 2.270 ;
        RECT  7.270 1.360 7.500 3.190 ;
        RECT  7.080 1.360 7.270 1.700 ;
        RECT  7.160 2.850 7.270 3.190 ;
        RECT  5.590 2.905 7.160 3.135 ;
        RECT  5.525 0.875 5.755 1.775 ;
        RECT  5.360 2.220 5.590 3.135 ;
        RECT  5.015 1.545 5.525 1.775 ;
        RECT  5.250 2.220 5.360 2.560 ;
        RECT  4.785 1.545 5.015 2.985 ;
        RECT  4.560 0.960 4.900 1.300 ;
        RECT  4.560 3.260 4.900 3.710 ;
        RECT  2.665 2.755 4.785 2.985 ;
        RECT  3.430 1.070 4.560 1.300 ;
        RECT  1.780 3.260 4.560 3.490 ;
        RECT  3.200 1.070 3.430 1.440 ;
        RECT  1.880 1.210 3.200 1.440 ;
        RECT  2.435 2.320 2.665 2.985 ;
        RECT  2.150 2.320 2.435 2.550 ;
        RECT  1.810 2.210 2.150 2.550 ;
        RECT  1.580 1.210 1.880 1.550 ;
        RECT  1.580 3.060 1.780 3.870 ;
        RECT  1.440 1.210 1.580 3.870 ;
        RECT  1.350 1.210 1.440 3.600 ;
        RECT  1.080 0.720 1.270 0.950 ;
        RECT  0.850 0.720 1.080 3.735 ;
        RECT  0.740 1.275 0.850 1.615 ;
        RECT  0.740 2.925 0.850 3.735 ;
    END
END TLATNSRX2

MACRO TLATNSRX1
    CLASS CORE ;
    FOREIGN TLATNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSRXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.105 0.555 2.445 ;
        RECT  0.140 1.840 0.545 2.445 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 2.130 3.850 2.470 ;
        RECT  3.510 1.845 3.820 2.470 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 1.310 11.040 3.360 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.640 2.965 9.685 3.205 ;
        RECT  9.620 2.965 9.640 3.310 ;
        RECT  9.390 1.430 9.620 3.310 ;
        RECT  9.280 1.430 9.390 1.770 ;
        RECT  9.300 2.970 9.390 3.310 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 1.930 6.900 2.270 ;
        RECT  6.385 1.930 6.560 2.160 ;
        RECT  6.155 1.845 6.385 2.160 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.900 3.085 2.660 ;
        RECT  2.580 1.900 2.780 2.240 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 -0.400 11.220 0.400 ;
        RECT  9.980 -0.400 10.320 0.575 ;
        RECT  8.820 -0.400 9.980 0.400 ;
        RECT  8.480 -0.400 8.820 0.575 ;
        RECT  6.710 -0.400 8.480 0.400 ;
        RECT  6.370 -0.400 6.710 0.575 ;
        RECT  2.720 -0.400 6.370 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  0.520 -0.400 2.380 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.375 4.640 11.220 5.440 ;
        RECT  9.975 4.465 10.375 5.440 ;
        RECT  8.880 4.640 9.975 5.440 ;
        RECT  8.540 4.465 8.880 5.440 ;
        RECT  6.820 4.640 8.540 5.440 ;
        RECT  6.480 4.465 6.820 5.440 ;
        RECT  3.500 4.640 6.480 5.440 ;
        RECT  3.160 4.135 3.500 5.440 ;
        RECT  0.520 4.640 3.160 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.415 2.070 10.470 2.410 ;
        RECT  10.185 0.805 10.415 4.015 ;
        RECT  9.620 0.805 10.185 1.035 ;
        RECT  10.130 2.070 10.185 2.410 ;
        RECT  9.640 3.785 10.185 4.015 ;
        RECT  9.410 3.785 9.640 4.365 ;
        RECT  9.280 0.635 9.620 1.035 ;
        RECT  9.300 4.005 9.410 4.365 ;
        RECT  5.950 4.005 9.300 4.235 ;
        RECT  9.025 2.090 9.160 2.430 ;
        RECT  8.795 2.090 9.025 3.775 ;
        RECT  4.820 3.545 8.795 3.775 ;
        RECT  7.965 0.765 8.195 3.170 ;
        RECT  7.680 0.765 7.965 1.105 ;
        RECT  7.780 2.830 7.965 3.170 ;
        RECT  7.485 1.900 7.730 2.240 ;
        RECT  5.655 0.875 7.680 1.105 ;
        RECT  7.255 1.365 7.485 3.315 ;
        RECT  6.980 1.365 7.255 1.595 ;
        RECT  7.075 2.570 7.255 3.315 ;
        RECT  5.190 2.570 7.075 2.800 ;
        RECT  5.425 0.875 5.655 1.940 ;
        RECT  5.010 1.710 5.425 1.940 ;
        RECT  4.850 2.460 5.190 2.800 ;
        RECT  4.670 1.710 5.010 2.050 ;
        RECT  4.480 3.370 4.820 3.775 ;
        RECT  4.450 1.820 4.670 2.050 ;
        RECT  4.260 1.040 4.600 1.380 ;
        RECT  1.820 3.545 4.480 3.775 ;
        RECT  4.220 1.820 4.450 3.135 ;
        RECT  2.595 1.150 4.260 1.380 ;
        RECT  2.475 2.905 4.220 3.135 ;
        RECT  2.365 1.150 2.595 1.545 ;
        RECT  2.245 2.470 2.475 3.135 ;
        RECT  1.620 1.315 2.365 1.545 ;
        RECT  2.190 2.470 2.245 2.700 ;
        RECT  1.850 2.360 2.190 2.700 ;
        RECT  1.620 0.730 1.960 1.070 ;
        RECT  1.620 3.110 1.820 3.775 ;
        RECT  1.290 4.020 1.630 4.360 ;
        RECT  1.120 0.840 1.620 1.070 ;
        RECT  1.590 1.315 1.620 3.775 ;
        RECT  1.390 1.315 1.590 3.450 ;
        RECT  1.120 4.020 1.290 4.250 ;
        RECT  0.890 0.840 1.120 4.250 ;
        RECT  0.780 1.290 0.890 1.630 ;
        RECT  0.780 2.930 0.890 3.270 ;
    END
END TLATNSRX1

MACRO TLATNSXL
    CLASS CORE ;
    FOREIGN TLATNSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 2.015 0.560 2.355 ;
        RECT  0.140 1.820 0.550 2.355 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 1.270 10.360 1.845 ;
        RECT  10.345 3.020 10.360 3.360 ;
        RECT  10.115 1.270 10.345 3.360 ;
        RECT  10.040 1.270 10.115 1.845 ;
        RECT  10.020 3.020 10.115 3.360 ;
        RECT  10.020 1.270 10.040 1.610 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.925 1.400 9.155 3.310 ;
        RECT  8.640 1.400 8.925 1.740 ;
        RECT  8.680 2.940 8.925 3.310 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.890 1.500 6.230 1.840 ;
        RECT  5.725 1.500 5.890 1.730 ;
        RECT  5.495 1.285 5.725 1.730 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.845 3.440 2.185 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.720 -0.400 10.560 0.400 ;
        RECT  9.380 -0.400 9.720 0.575 ;
        RECT  8.170 -0.400 9.380 0.400 ;
        RECT  7.830 -0.400 8.170 0.575 ;
        RECT  5.770 -0.400 7.830 0.400 ;
        RECT  5.430 -0.400 5.770 0.575 ;
        RECT  2.740 -0.400 5.430 0.400 ;
        RECT  2.400 -0.400 2.740 0.575 ;
        RECT  0.520 -0.400 2.400 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.765 4.640 10.560 5.440 ;
        RECT  9.355 4.465 9.765 5.440 ;
        RECT  8.260 4.640 9.355 5.440 ;
        RECT  7.920 4.465 8.260 5.440 ;
        RECT  6.200 4.640 7.920 5.440 ;
        RECT  5.860 4.465 6.200 5.440 ;
        RECT  3.460 4.640 5.860 5.440 ;
        RECT  3.120 4.005 3.460 5.440 ;
        RECT  0.520 4.640 3.120 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.630 2.070 9.740 2.410 ;
        RECT  9.400 0.885 9.630 4.015 ;
        RECT  9.125 0.885 9.400 1.115 ;
        RECT  9.040 3.785 9.400 4.015 ;
        RECT  8.895 0.665 9.125 1.115 ;
        RECT  8.810 3.785 9.040 4.365 ;
        RECT  8.680 0.665 8.895 0.895 ;
        RECT  8.680 4.005 8.810 4.365 ;
        RECT  5.330 4.005 8.680 4.235 ;
        RECT  8.205 2.070 8.540 2.410 ;
        RECT  7.975 2.070 8.205 3.775 ;
        RECT  1.780 3.545 7.975 3.775 ;
        RECT  7.270 1.290 7.500 3.315 ;
        RECT  7.010 1.290 7.270 1.630 ;
        RECT  7.160 2.885 7.270 3.315 ;
        RECT  4.015 3.085 7.160 3.315 ;
        RECT  6.825 1.935 7.035 2.290 ;
        RECT  6.695 1.935 6.825 2.855 ;
        RECT  6.465 0.850 6.695 2.855 ;
        RECT  6.270 0.850 6.465 1.190 ;
        RECT  4.680 2.625 6.465 2.855 ;
        RECT  4.450 2.260 4.680 2.855 ;
        RECT  4.330 1.500 4.670 1.840 ;
        RECT  4.340 2.260 4.450 2.600 ;
        RECT  4.050 0.830 4.390 1.170 ;
        RECT  4.015 1.610 4.330 1.840 ;
        RECT  3.315 0.940 4.050 1.170 ;
        RECT  3.785 1.610 4.015 3.315 ;
        RECT  2.095 2.495 3.785 2.725 ;
        RECT  3.085 0.940 3.315 1.565 ;
        RECT  1.585 1.335 3.085 1.565 ;
        RECT  1.865 2.360 2.095 2.725 ;
        RECT  1.120 0.765 1.930 0.995 ;
        RECT  1.585 3.110 1.780 3.775 ;
        RECT  1.250 4.020 1.590 4.360 ;
        RECT  1.495 1.335 1.585 3.775 ;
        RECT  1.355 1.335 1.495 3.450 ;
        RECT  1.120 4.020 1.250 4.250 ;
        RECT  0.890 0.765 1.120 4.250 ;
        RECT  0.780 1.330 0.890 1.670 ;
        RECT  0.740 2.980 0.890 3.320 ;
    END
END TLATNSXL

MACRO TLATNSX4
    CLASS CORE ;
    FOREIGN TLATNSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.090 0.555 2.430 ;
        RECT  0.140 1.845 0.545 2.430 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.040 1.515 13.060 3.220 ;
        RECT  12.700 1.360 13.040 3.220 ;
        RECT  12.680 1.515 12.700 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.740 1.360 11.760 1.940 ;
        RECT  11.740 2.880 11.760 3.220 ;
        RECT  11.420 1.360 11.740 3.220 ;
        RECT  11.360 1.820 11.420 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  7.780 1.420 7.865 1.770 ;
        RECT  7.475 1.420 7.780 2.100 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.250 2.070 3.360 2.580 ;
        RECT  3.020 1.845 3.250 2.580 ;
        RECT  2.855 1.845 3.020 2.075 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.680 -0.400 13.860 0.400 ;
        RECT  13.340 -0.400 13.680 0.950 ;
        RECT  12.400 -0.400 13.340 0.400 ;
        RECT  12.060 -0.400 12.400 0.950 ;
        RECT  11.120 -0.400 12.060 0.400 ;
        RECT  10.780 -0.400 11.120 0.950 ;
        RECT  9.700 -0.400 10.780 0.400 ;
        RECT  9.360 -0.400 9.700 1.305 ;
        RECT  7.480 -0.400 9.360 0.400 ;
        RECT  7.140 -0.400 7.480 0.575 ;
        RECT  5.400 -0.400 7.140 0.400 ;
        RECT  5.060 -0.400 5.400 0.575 ;
        RECT  2.700 -0.400 5.060 0.400 ;
        RECT  2.360 -0.400 2.700 0.575 ;
        RECT  0.520 -0.400 2.360 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.680 4.640 13.860 5.440 ;
        RECT  13.340 4.090 13.680 5.440 ;
        RECT  12.400 4.640 13.340 5.440 ;
        RECT  12.060 4.090 12.400 5.440 ;
        RECT  11.080 4.640 12.060 5.440 ;
        RECT  10.740 4.465 11.080 5.440 ;
        RECT  9.840 4.640 10.740 5.440 ;
        RECT  9.500 4.465 9.840 5.440 ;
        RECT  8.020 4.640 9.500 5.440 ;
        RECT  7.680 4.465 8.020 5.440 ;
        RECT  3.620 4.640 7.680 5.440 ;
        RECT  3.280 3.815 3.620 5.440 ;
        RECT  0.520 4.640 3.280 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 2.070 13.670 2.410 ;
        RECT  13.385 2.070 13.615 3.810 ;
        RECT  13.330 2.070 13.385 2.410 ;
        RECT  10.500 3.580 13.385 3.810 ;
        RECT  10.880 1.330 11.110 3.060 ;
        RECT  10.420 1.330 10.880 1.560 ;
        RECT  10.500 2.830 10.880 3.060 ;
        RECT  9.865 2.070 10.650 2.410 ;
        RECT  10.445 2.830 10.500 4.175 ;
        RECT  10.160 2.830 10.445 4.195 ;
        RECT  10.080 1.220 10.420 1.560 ;
        RECT  7.150 3.965 10.160 4.195 ;
        RECT  9.635 2.070 9.865 3.635 ;
        RECT  5.670 3.405 9.635 3.635 ;
        RECT  9.065 2.945 9.180 3.175 ;
        RECT  8.835 0.955 9.065 3.175 ;
        RECT  8.600 0.955 8.835 1.295 ;
        RECT  5.975 2.945 8.835 3.175 ;
        RECT  8.480 1.605 8.535 1.975 ;
        RECT  8.325 1.605 8.480 2.625 ;
        RECT  8.095 0.810 8.325 2.625 ;
        RECT  7.900 0.810 8.095 1.150 ;
        RECT  6.630 2.395 8.095 2.625 ;
        RECT  6.265 2.275 6.630 2.625 ;
        RECT  6.070 1.400 6.410 1.740 ;
        RECT  5.780 0.830 6.120 1.170 ;
        RECT  5.975 1.510 6.070 1.740 ;
        RECT  5.745 1.510 5.975 3.175 ;
        RECT  5.225 0.940 5.780 1.170 ;
        RECT  5.490 2.600 5.745 2.940 ;
        RECT  5.330 3.405 5.670 3.770 ;
        RECT  4.245 2.710 5.490 2.940 ;
        RECT  4.675 3.405 5.330 3.635 ;
        RECT  4.995 0.940 5.225 1.190 ;
        RECT  4.050 0.960 4.995 1.190 ;
        RECT  4.445 3.355 4.675 3.635 ;
        RECT  1.780 3.355 4.445 3.585 ;
        RECT  4.015 2.710 4.245 3.120 ;
        RECT  3.995 0.960 4.050 1.300 ;
        RECT  2.250 2.890 4.015 3.120 ;
        RECT  3.710 0.960 3.995 1.480 ;
        RECT  1.780 1.250 3.710 1.480 ;
        RECT  2.020 2.235 2.250 3.120 ;
        RECT  1.825 2.235 2.020 2.580 ;
        RECT  1.080 0.765 1.930 0.995 ;
        RECT  1.770 2.240 1.825 2.580 ;
        RECT  1.540 1.250 1.780 1.590 ;
        RECT  1.540 3.320 1.780 3.660 ;
        RECT  1.310 1.250 1.540 3.660 ;
        RECT  0.850 0.765 1.080 3.540 ;
        RECT  0.740 1.250 0.850 1.590 ;
        RECT  0.740 3.200 0.850 3.540 ;
    END
END TLATNSX4

MACRO TLATNSX2
    CLASS CORE ;
    FOREIGN TLATNSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 2.080 0.555 2.420 ;
        RECT  0.140 1.840 0.545 2.420 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.025 2.940 11.040 4.220 ;
        RECT  10.700 0.835 11.025 4.220 ;
        RECT  10.685 0.835 10.700 3.750 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.765 1.335 9.995 3.050 ;
        RECT  9.060 1.335 9.765 1.565 ;
        RECT  9.600 2.820 9.765 3.050 ;
        RECT  9.260 2.820 9.600 3.195 ;
        RECT  8.795 2.910 9.260 3.195 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 1.500 6.130 1.840 ;
        RECT  5.725 1.500 5.790 1.730 ;
        RECT  5.495 1.285 5.725 1.730 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.845 3.390 2.185 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.220 -0.400 11.220 0.400 ;
        RECT  9.880 -0.400 10.220 0.575 ;
        RECT  7.960 -0.400 9.880 0.400 ;
        RECT  7.620 -0.400 7.960 1.585 ;
        RECT  5.660 -0.400 7.620 0.400 ;
        RECT  5.320 -0.400 5.660 0.575 ;
        RECT  2.880 -0.400 5.320 0.400 ;
        RECT  2.540 -0.400 2.880 0.575 ;
        RECT  0.520 -0.400 2.540 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 4.640 11.220 5.440 ;
        RECT  9.980 4.080 10.320 5.440 ;
        RECT  8.200 4.640 9.980 5.440 ;
        RECT  7.860 4.465 8.200 5.440 ;
        RECT  6.200 4.640 7.860 5.440 ;
        RECT  5.860 4.465 6.200 5.440 ;
        RECT  3.700 4.640 5.860 5.440 ;
        RECT  3.360 4.090 3.700 5.440 ;
        RECT  0.520 4.640 3.360 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.225 0.870 10.455 3.850 ;
        RECT  8.680 0.870 10.225 1.100 ;
        RECT  8.960 3.620 10.225 3.850 ;
        RECT  8.205 2.070 9.060 2.410 ;
        RECT  8.850 3.620 8.960 3.960 ;
        RECT  8.620 3.620 8.850 4.225 ;
        RECT  8.450 0.870 8.680 1.585 ;
        RECT  5.330 3.995 8.620 4.225 ;
        RECT  8.340 1.245 8.450 1.585 ;
        RECT  7.975 2.070 8.205 3.735 ;
        RECT  4.200 3.505 7.975 3.735 ;
        RECT  7.390 2.855 7.500 3.275 ;
        RECT  7.160 1.245 7.390 3.275 ;
        RECT  6.820 1.245 7.160 1.585 ;
        RECT  4.790 3.045 7.160 3.275 ;
        RECT  6.825 1.890 6.915 2.275 ;
        RECT  6.590 1.890 6.825 2.815 ;
        RECT  6.360 0.850 6.590 2.815 ;
        RECT  6.120 0.850 6.360 1.190 ;
        RECT  5.255 2.585 6.360 2.815 ;
        RECT  5.025 2.505 5.255 2.815 ;
        RECT  4.230 2.505 5.025 2.735 ;
        RECT  4.560 2.965 4.790 3.275 ;
        RECT  4.310 1.780 4.650 2.120 ;
        RECT  3.925 2.965 4.560 3.195 ;
        RECT  3.925 1.890 4.310 2.120 ;
        RECT  3.960 0.810 4.300 1.150 ;
        RECT  3.860 3.425 4.200 3.735 ;
        RECT  2.475 0.865 3.960 1.095 ;
        RECT  3.695 1.890 3.925 3.195 ;
        RECT  1.820 3.505 3.860 3.735 ;
        RECT  2.475 2.965 3.695 3.195 ;
        RECT  2.245 0.865 2.475 1.490 ;
        RECT  2.245 2.230 2.475 3.195 ;
        RECT  1.900 1.260 2.245 1.490 ;
        RECT  2.190 2.230 2.245 2.460 ;
        RECT  1.850 2.120 2.190 2.460 ;
        RECT  1.120 0.765 1.930 0.995 ;
        RECT  1.620 1.260 1.900 1.600 ;
        RECT  1.620 2.775 1.820 4.055 ;
        RECT  1.480 1.260 1.620 4.055 ;
        RECT  1.390 1.260 1.480 3.735 ;
        RECT  0.890 0.765 1.120 3.120 ;
        RECT  0.780 1.290 0.890 1.630 ;
        RECT  0.780 2.780 0.890 3.120 ;
    END
END TLATNSX2

MACRO TLATNSX1
    CLASS CORE ;
    FOREIGN TLATNSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 2.015 0.560 2.355 ;
        RECT  0.140 1.820 0.550 2.355 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 1.320 10.360 1.845 ;
        RECT  10.345 3.020 10.360 3.360 ;
        RECT  10.115 1.320 10.345 3.360 ;
        RECT  10.040 1.320 10.115 1.845 ;
        RECT  10.020 3.020 10.115 3.360 ;
        RECT  10.020 1.320 10.040 1.770 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.135 1.430 9.155 3.195 ;
        RECT  8.925 1.430 9.135 3.310 ;
        RECT  8.660 1.430 8.925 1.770 ;
        RECT  8.680 2.940 8.925 3.310 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.890 1.500 6.230 1.840 ;
        RECT  5.725 1.500 5.890 1.730 ;
        RECT  5.495 1.285 5.725 1.730 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 1.845 3.460 2.185 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.720 -0.400 10.560 0.400 ;
        RECT  9.380 -0.400 9.720 0.575 ;
        RECT  8.170 -0.400 9.380 0.400 ;
        RECT  7.830 -0.400 8.170 0.575 ;
        RECT  5.770 -0.400 7.830 0.400 ;
        RECT  5.430 -0.400 5.770 0.575 ;
        RECT  2.740 -0.400 5.430 0.400 ;
        RECT  2.400 -0.400 2.740 0.575 ;
        RECT  0.520 -0.400 2.400 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.775 4.640 10.560 5.440 ;
        RECT  9.355 4.465 9.775 5.440 ;
        RECT  8.260 4.640 9.355 5.440 ;
        RECT  7.920 4.465 8.260 5.440 ;
        RECT  6.200 4.640 7.920 5.440 ;
        RECT  5.860 4.465 6.200 5.440 ;
        RECT  3.460 4.640 5.860 5.440 ;
        RECT  3.120 4.110 3.460 5.440 ;
        RECT  0.520 4.640 3.120 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.630 2.070 9.740 2.410 ;
        RECT  9.400 0.885 9.630 4.015 ;
        RECT  9.125 0.885 9.400 1.115 ;
        RECT  9.020 3.785 9.400 4.015 ;
        RECT  8.895 0.655 9.125 1.115 ;
        RECT  8.790 3.785 9.020 4.365 ;
        RECT  8.680 0.655 8.895 0.885 ;
        RECT  8.680 4.005 8.790 4.365 ;
        RECT  5.330 4.005 8.680 4.235 ;
        RECT  8.205 2.070 8.540 2.410 ;
        RECT  7.975 2.070 8.205 3.775 ;
        RECT  1.780 3.545 7.975 3.775 ;
        RECT  7.270 0.650 7.500 3.315 ;
        RECT  6.990 0.650 7.270 0.990 ;
        RECT  7.160 2.885 7.270 3.315 ;
        RECT  4.015 3.085 7.160 3.315 ;
        RECT  6.825 1.635 7.035 2.015 ;
        RECT  6.695 1.635 6.825 2.855 ;
        RECT  6.465 0.850 6.695 2.855 ;
        RECT  6.270 0.850 6.465 1.190 ;
        RECT  4.680 2.625 6.465 2.855 ;
        RECT  4.450 2.260 4.680 2.855 ;
        RECT  4.330 1.500 4.670 1.840 ;
        RECT  4.340 2.260 4.450 2.600 ;
        RECT  4.030 0.810 4.370 1.150 ;
        RECT  4.015 1.610 4.330 1.840 ;
        RECT  3.315 0.920 4.030 1.150 ;
        RECT  3.785 1.610 4.015 3.315 ;
        RECT  2.095 2.495 3.785 2.725 ;
        RECT  3.085 0.920 3.315 1.565 ;
        RECT  1.900 1.335 3.085 1.565 ;
        RECT  1.865 2.360 2.095 2.725 ;
        RECT  1.590 0.700 1.930 1.040 ;
        RECT  1.585 1.280 1.900 1.620 ;
        RECT  1.585 3.110 1.780 3.775 ;
        RECT  1.120 0.810 1.590 1.040 ;
        RECT  1.250 4.020 1.590 4.360 ;
        RECT  1.560 1.280 1.585 3.775 ;
        RECT  1.495 1.335 1.560 3.775 ;
        RECT  1.355 1.335 1.495 3.450 ;
        RECT  1.120 4.020 1.250 4.250 ;
        RECT  0.890 0.810 1.120 4.250 ;
        RECT  0.780 1.330 0.890 1.670 ;
        RECT  0.740 2.980 0.890 3.320 ;
    END
END TLATNSX1

MACRO TLATNRXL
    CLASS CORE ;
    FOREIGN TLATNRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 2.405 5.065 2.635 ;
        RECT  4.740 2.060 4.850 2.660 ;
        RECT  4.510 2.060 4.740 2.885 ;
        RECT  3.745 2.655 4.510 2.885 ;
        RECT  3.405 2.655 3.745 3.130 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 1.230 8.400 3.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.505 0.810 7.735 3.755 ;
        RECT  6.960 0.810 7.505 1.040 ;
        RECT  7.140 3.525 7.505 3.755 ;
        RECT  6.815 3.525 7.140 4.015 ;
        RECT  6.620 0.700 6.960 1.040 ;
        RECT  6.800 3.555 6.815 4.015 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.530 2.520 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.405 2.425 3.150 ;
        RECT  1.995 2.810 2.120 3.150 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.720 -0.400 8.580 0.400 ;
        RECT  7.380 -0.400 7.720 0.575 ;
        RECT  6.080 -0.400 7.380 0.400 ;
        RECT  5.740 -0.400 6.080 0.575 ;
        RECT  2.020 -0.400 5.740 0.400 ;
        RECT  1.680 -0.400 2.020 0.575 ;
        RECT  0.520 -0.400 1.680 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.780 4.640 8.580 5.440 ;
        RECT  7.375 4.465 7.780 5.440 ;
        RECT  6.380 4.640 7.375 5.440 ;
        RECT  6.040 4.465 6.380 5.440 ;
        RECT  4.175 4.640 6.040 5.440 ;
        RECT  3.835 3.850 4.175 5.440 ;
        RECT  2.095 4.640 3.835 5.440 ;
        RECT  1.755 3.570 2.095 5.440 ;
        RECT  0.520 4.640 1.755 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.045 1.565 7.275 3.175 ;
        RECT  6.960 1.565 7.045 1.795 ;
        RECT  6.800 2.810 7.045 3.175 ;
        RECT  6.620 1.455 6.960 1.795 ;
        RECT  6.395 2.945 6.800 3.175 ;
        RECT  6.320 2.070 6.660 2.410 ;
        RECT  6.165 2.945 6.395 4.070 ;
        RECT  5.835 2.125 6.320 2.355 ;
        RECT  5.820 3.840 6.165 4.070 ;
        RECT  5.825 2.125 5.835 3.460 ;
        RECT  5.605 1.170 5.825 3.460 ;
        RECT  5.480 3.840 5.820 4.180 ;
        RECT  5.595 1.170 5.605 2.355 ;
        RECT  4.935 3.230 5.605 3.460 ;
        RECT  3.900 1.170 5.595 1.400 ;
        RECT  4.570 3.230 4.935 3.620 ;
        RECT  3.375 3.390 4.570 3.620 ;
        RECT  3.840 1.630 4.180 1.970 ;
        RECT  3.560 1.060 3.900 1.400 ;
        RECT  3.015 1.685 3.840 1.915 ;
        RECT  3.035 3.390 3.375 3.770 ;
        RECT  3.015 2.790 3.070 3.130 ;
        RECT  2.785 1.685 3.015 3.130 ;
        RECT  1.675 1.685 2.785 1.915 ;
        RECT  2.730 2.790 2.785 3.130 ;
        RECT  1.525 0.805 1.675 3.175 ;
        RECT  1.445 0.805 1.525 3.910 ;
        RECT  1.220 0.805 1.445 1.040 ;
        RECT  1.295 2.945 1.445 3.910 ;
        RECT  1.035 3.570 1.295 3.910 ;
        RECT  0.880 0.700 1.220 1.040 ;
        RECT  1.065 2.270 1.215 2.610 ;
        RECT  1.065 1.400 1.120 1.740 ;
        RECT  0.835 1.400 1.065 3.190 ;
        RECT  0.780 1.400 0.835 1.740 ;
    END
END TLATNRXL

MACRO TLATNRX4
    CLASS CORE ;
    FOREIGN TLATNRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.600 3.400 2.940 ;
        RECT  2.855 2.405 3.085 2.940 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.060 1.820 11.080 3.220 ;
        RECT  10.720 1.455 11.060 3.220 ;
        RECT  10.700 1.820 10.720 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.760 1.455 9.780 1.845 ;
        RECT  9.760 2.635 9.780 3.180 ;
        RECT  9.440 1.455 9.760 3.220 ;
        RECT  9.380 1.820 9.440 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  5.715 1.750 6.295 2.100 ;
        RECT  5.495 1.845 5.715 2.075 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 1.845 1.990 2.340 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.700 -0.400 11.880 0.400 ;
        RECT  11.360 -0.400 11.700 1.045 ;
        RECT  10.420 -0.400 11.360 0.400 ;
        RECT  10.080 -0.400 10.420 1.045 ;
        RECT  9.100 -0.400 10.080 0.400 ;
        RECT  8.760 -0.400 9.100 0.575 ;
        RECT  7.200 -0.400 8.760 0.400 ;
        RECT  6.160 -0.400 7.200 0.575 ;
        RECT  2.440 -0.400 6.160 0.400 ;
        RECT  2.100 -0.400 2.440 1.055 ;
        RECT  0.000 -0.400 2.100 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.700 4.640 11.880 5.440 ;
        RECT  11.360 4.090 11.700 5.440 ;
        RECT  10.420 4.640 11.360 5.440 ;
        RECT  10.080 4.090 10.420 5.440 ;
        RECT  9.140 4.640 10.080 5.440 ;
        RECT  8.800 4.090 9.140 5.440 ;
        RECT  7.620 4.640 8.800 5.440 ;
        RECT  7.280 4.465 7.620 5.440 ;
        RECT  5.360 4.640 7.280 5.440 ;
        RECT  5.020 4.465 5.360 5.440 ;
        RECT  3.120 4.640 5.020 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  0.520 4.640 2.780 5.440 ;
        RECT  0.180 4.145 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.615 2.100 11.670 2.440 ;
        RECT  11.385 2.100 11.615 3.860 ;
        RECT  11.330 2.100 11.385 2.440 ;
        RECT  8.865 3.630 11.385 3.860 ;
        RECT  8.635 1.565 8.865 3.860 ;
        RECT  8.500 1.565 8.635 1.795 ;
        RECT  8.345 3.570 8.635 3.860 ;
        RECT  8.160 1.455 8.500 1.795 ;
        RECT  8.115 3.570 8.345 4.175 ;
        RECT  8.230 2.200 8.340 2.540 ;
        RECT  8.000 2.200 8.230 3.340 ;
        RECT  4.775 3.945 8.115 4.175 ;
        RECT  7.885 3.110 8.000 3.340 ;
        RECT  7.960 0.705 7.965 1.095 ;
        RECT  7.770 0.650 7.960 1.095 ;
        RECT  7.655 3.110 7.885 3.655 ;
        RECT  7.620 0.650 7.770 2.875 ;
        RECT  3.920 3.425 7.655 3.655 ;
        RECT  7.540 0.865 7.620 2.875 ;
        RECT  4.785 0.865 7.540 1.095 ;
        RECT  7.425 2.645 7.540 2.875 ;
        RECT  7.195 2.645 7.425 3.080 ;
        RECT  6.965 1.955 7.245 2.320 ;
        RECT  6.860 2.850 7.195 3.080 ;
        RECT  6.735 1.410 6.965 2.615 ;
        RECT  6.520 2.850 6.860 3.190 ;
        RECT  6.615 1.410 6.735 1.750 ;
        RECT  6.160 2.385 6.735 2.615 ;
        RECT  5.930 2.385 6.160 3.190 ;
        RECT  5.820 2.850 5.930 3.190 ;
        RECT  4.675 2.850 5.820 3.080 ;
        RECT  4.555 0.865 4.785 2.260 ;
        RECT  4.545 3.945 4.775 4.310 ;
        RECT  4.445 2.765 4.675 3.080 ;
        RECT  4.350 1.875 4.555 2.260 ;
        RECT  4.080 2.765 4.445 2.995 ;
        RECT  2.475 1.875 4.350 2.105 ;
        RECT  4.265 0.980 4.320 1.320 ;
        RECT  3.980 0.980 4.265 1.515 ;
        RECT  3.820 3.970 4.160 4.310 ;
        RECT  3.795 2.650 4.080 2.995 ;
        RECT  1.035 1.285 3.980 1.515 ;
        RECT  3.580 3.290 3.920 3.655 ;
        RECT  2.355 3.970 3.820 4.200 ;
        RECT  3.740 2.650 3.795 2.990 ;
        RECT  1.800 3.425 3.580 3.655 ;
        RECT  2.245 1.875 2.475 2.955 ;
        RECT  2.125 3.970 2.355 4.285 ;
        RECT  1.460 2.725 2.245 2.955 ;
        RECT  1.125 4.055 2.125 4.285 ;
        RECT  1.690 3.425 1.800 3.820 ;
        RECT  1.460 3.220 1.690 3.820 ;
        RECT  1.035 3.220 1.460 3.450 ;
        RECT  0.895 3.685 1.125 4.285 ;
        RECT  0.805 1.285 1.035 3.450 ;
        RECT  0.495 3.685 0.895 3.915 ;
        RECT  0.520 1.285 0.805 1.515 ;
        RECT  0.180 1.120 0.520 1.515 ;
        RECT  0.265 1.820 0.495 3.915 ;
    END
END TLATNRX4

MACRO TLATNRX2
    CLASS CORE ;
    FOREIGN TLATNRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNRXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 2.940 4.450 3.220 ;
        RECT  4.300 2.940 4.410 3.510 ;
        RECT  4.070 2.275 4.300 3.510 ;
        RECT  3.390 2.275 4.070 2.505 ;
        RECT  3.160 1.895 3.390 2.505 ;
        RECT  3.050 1.895 3.160 2.125 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.025 0.765 9.060 1.575 ;
        RECT  9.025 2.970 9.060 4.250 ;
        RECT  8.795 0.765 9.025 4.250 ;
        RECT  8.720 0.765 8.795 1.575 ;
        RECT  8.720 2.970 8.795 4.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.540 2.965 7.705 3.195 ;
        RECT  7.485 1.390 7.540 1.845 ;
        RECT  7.485 2.965 7.540 4.250 ;
        RECT  7.255 1.390 7.485 4.250 ;
        RECT  7.200 1.390 7.255 1.730 ;
        RECT  7.200 2.970 7.255 4.250 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.530 2.575 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 2.190 2.700 2.660 ;
        RECT  2.025 2.230 2.360 2.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 -0.400 9.240 0.400 ;
        RECT  7.960 -0.400 8.300 0.575 ;
        RECT  6.080 -0.400 7.960 0.400 ;
        RECT  5.740 -0.400 6.080 0.575 ;
        RECT  2.420 -0.400 5.740 0.400 ;
        RECT  2.080 -0.400 2.420 0.575 ;
        RECT  0.520 -0.400 2.080 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 4.640 9.240 5.440 ;
        RECT  7.960 4.465 8.300 5.440 ;
        RECT  6.270 4.640 7.960 5.440 ;
        RECT  5.855 4.465 6.270 5.440 ;
        RECT  4.200 4.640 5.855 5.440 ;
        RECT  3.860 4.465 4.200 5.440 ;
        RECT  2.120 4.640 3.860 5.440 ;
        RECT  1.780 4.090 2.120 5.440 ;
        RECT  0.520 4.640 1.780 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.340 2.100 8.450 2.440 ;
        RECT  8.110 0.865 8.340 2.440 ;
        RECT  6.840 0.865 8.110 1.095 ;
        RECT  6.785 0.640 6.840 1.095 ;
        RECT  6.785 3.020 6.840 3.360 ;
        RECT  6.555 0.640 6.785 3.360 ;
        RECT  6.500 0.640 6.555 0.980 ;
        RECT  6.060 1.620 6.555 1.960 ;
        RECT  6.500 3.020 6.555 3.360 ;
        RECT  5.725 2.315 6.315 2.705 ;
        RECT  5.495 0.890 5.725 4.135 ;
        RECT  4.300 0.890 5.495 1.120 ;
        RECT  3.400 3.905 5.495 4.135 ;
        RECT  5.070 3.295 5.180 3.635 ;
        RECT  4.840 1.815 5.070 3.635 ;
        RECT  3.950 1.815 4.840 2.045 ;
        RECT  3.960 0.780 4.300 1.120 ;
        RECT  3.720 1.435 3.950 2.045 ;
        RECT  2.525 1.435 3.720 1.665 ;
        RECT  3.060 3.905 3.400 4.350 ;
        RECT  3.210 2.735 3.370 2.965 ;
        RECT  2.980 2.735 3.210 3.245 ;
        RECT  1.675 3.015 2.980 3.245 ;
        RECT  2.295 0.820 2.525 1.665 ;
        RECT  1.120 0.820 2.295 1.050 ;
        RECT  1.675 1.295 1.820 1.525 ;
        RECT  1.445 1.295 1.675 3.860 ;
        RECT  1.300 3.630 1.445 3.860 ;
        RECT  0.960 3.630 1.300 3.970 ;
        RECT  1.120 2.060 1.215 2.405 ;
        RECT  0.890 0.820 1.120 3.120 ;
        RECT  0.780 1.240 0.890 1.580 ;
        RECT  0.780 2.780 0.890 3.120 ;
    END
END TLATNRX2

MACRO TLATNRX1
    CLASS CORE ;
    FOREIGN TLATNRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNRXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 2.405 5.065 2.635 ;
        RECT  4.740 2.060 4.850 2.660 ;
        RECT  4.510 2.060 4.740 2.885 ;
        RECT  3.745 2.655 4.510 2.885 ;
        RECT  3.405 2.655 3.745 3.130 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 1.200 8.400 3.300 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.505 0.865 7.735 3.755 ;
        RECT  6.960 0.865 7.505 1.095 ;
        RECT  7.140 3.525 7.505 3.755 ;
        RECT  6.800 3.525 7.140 4.140 ;
        RECT  6.620 0.700 6.960 1.095 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.845 0.530 2.570 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.405 2.425 3.170 ;
        RECT  1.995 2.830 2.120 3.170 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.720 -0.400 8.580 0.400 ;
        RECT  7.380 -0.400 7.720 0.575 ;
        RECT  6.080 -0.400 7.380 0.400 ;
        RECT  5.740 -0.400 6.080 0.575 ;
        RECT  2.020 -0.400 5.740 0.400 ;
        RECT  1.680 -0.400 2.020 0.575 ;
        RECT  0.520 -0.400 1.680 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.840 4.640 8.580 5.440 ;
        RECT  7.500 4.465 7.840 5.440 ;
        RECT  6.380 4.640 7.500 5.440 ;
        RECT  6.040 4.465 6.380 5.440 ;
        RECT  4.175 4.640 6.040 5.440 ;
        RECT  3.835 3.850 4.175 5.440 ;
        RECT  2.095 4.640 3.835 5.440 ;
        RECT  1.755 3.620 2.095 5.440 ;
        RECT  0.520 4.640 1.755 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.045 1.600 7.275 3.175 ;
        RECT  6.960 1.600 7.045 1.830 ;
        RECT  6.800 2.810 7.045 3.175 ;
        RECT  6.620 1.490 6.960 1.830 ;
        RECT  6.395 2.945 6.800 3.175 ;
        RECT  6.320 2.070 6.660 2.410 ;
        RECT  6.165 2.945 6.395 4.125 ;
        RECT  5.835 2.125 6.320 2.355 ;
        RECT  5.480 3.895 6.165 4.125 ;
        RECT  5.825 2.125 5.835 3.460 ;
        RECT  5.605 1.070 5.825 3.460 ;
        RECT  5.595 1.070 5.605 2.355 ;
        RECT  4.935 3.230 5.605 3.460 ;
        RECT  3.900 1.070 5.595 1.300 ;
        RECT  4.570 3.230 4.935 3.620 ;
        RECT  3.375 3.390 4.570 3.620 ;
        RECT  3.840 1.610 4.180 1.950 ;
        RECT  3.560 0.960 3.900 1.300 ;
        RECT  3.015 1.665 3.840 1.895 ;
        RECT  3.035 3.390 3.375 3.730 ;
        RECT  3.015 2.790 3.070 3.130 ;
        RECT  2.785 1.665 3.015 3.130 ;
        RECT  1.675 1.665 2.785 1.895 ;
        RECT  2.730 2.790 2.785 3.130 ;
        RECT  1.525 0.805 1.675 3.175 ;
        RECT  1.445 0.805 1.525 3.960 ;
        RECT  1.220 0.805 1.445 1.040 ;
        RECT  1.295 2.945 1.445 3.960 ;
        RECT  1.035 3.620 1.295 3.960 ;
        RECT  0.880 0.700 1.220 1.040 ;
        RECT  1.065 2.270 1.215 2.610 ;
        RECT  1.065 1.400 1.120 1.740 ;
        RECT  0.835 1.400 1.065 3.190 ;
        RECT  0.780 1.400 0.835 1.740 ;
    END
END TLATNRX1

MACRO TLATNXL
    CLASS CORE ;
    FOREIGN TLATNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 3.090 7.080 3.430 ;
        RECT  7.045 1.160 7.060 1.500 ;
        RECT  6.815 1.160 7.045 3.430 ;
        RECT  6.720 1.160 6.815 1.500 ;
        RECT  6.740 3.090 6.815 3.430 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.225 0.865 6.455 3.755 ;
        RECT  6.080 0.865 6.225 1.285 ;
        RECT  5.620 3.525 6.225 3.755 ;
        RECT  5.530 0.865 6.080 1.095 ;
        RECT  5.280 3.525 5.620 4.150 ;
        RECT  5.175 0.685 5.530 1.095 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.845 0.530 2.495 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 1.845 2.425 2.690 ;
        RECT  1.995 2.350 2.120 2.690 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.350 -0.400 7.260 0.400 ;
        RECT  6.010 -0.400 6.350 0.575 ;
        RECT  4.700 -0.400 6.010 0.400 ;
        RECT  4.360 -0.400 4.700 0.575 ;
        RECT  2.020 -0.400 4.360 0.400 ;
        RECT  1.680 -0.400 2.020 0.575 ;
        RECT  0.520 -0.400 1.680 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.375 4.640 7.260 5.440 ;
        RECT  5.960 4.465 6.375 5.440 ;
        RECT  4.860 4.640 5.960 5.440 ;
        RECT  4.520 4.465 4.860 5.440 ;
        RECT  2.095 4.640 4.520 5.440 ;
        RECT  1.755 3.460 2.095 5.440 ;
        RECT  0.520 4.640 1.755 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.700 2.100 5.810 2.440 ;
        RECT  5.470 1.400 5.700 3.190 ;
        RECT  5.190 1.400 5.470 1.740 ;
        RECT  5.280 2.850 5.470 3.190 ;
        RECT  4.855 2.960 5.280 3.190 ;
        RECT  4.800 2.070 5.140 2.410 ;
        RECT  4.625 2.960 4.855 3.850 ;
        RECT  4.185 2.070 4.800 2.300 ;
        RECT  4.325 3.620 4.625 3.850 ;
        RECT  3.985 3.620 4.325 3.960 ;
        RECT  3.955 0.805 4.185 3.285 ;
        RECT  3.340 0.805 3.955 1.035 ;
        RECT  3.375 3.055 3.955 3.285 ;
        RECT  3.305 1.280 3.645 1.620 ;
        RECT  3.140 3.055 3.375 3.590 ;
        RECT  3.000 0.680 3.340 1.035 ;
        RECT  3.135 1.360 3.305 1.620 ;
        RECT  3.035 3.250 3.140 3.590 ;
        RECT  2.905 1.360 3.135 2.765 ;
        RECT  1.675 1.360 2.905 1.590 ;
        RECT  2.795 2.535 2.905 2.765 ;
        RECT  1.525 0.865 1.675 3.135 ;
        RECT  1.445 0.865 1.525 3.690 ;
        RECT  1.220 0.865 1.445 1.095 ;
        RECT  1.295 2.905 1.445 3.690 ;
        RECT  1.260 3.460 1.295 3.690 ;
        RECT  0.920 3.460 1.260 3.800 ;
        RECT  0.880 0.805 1.220 1.095 ;
        RECT  1.120 2.060 1.215 2.405 ;
        RECT  1.065 1.450 1.120 2.405 ;
        RECT  0.890 1.450 1.065 3.080 ;
        RECT  0.780 1.450 0.890 1.790 ;
        RECT  0.835 2.175 0.890 3.080 ;
    END
END TLATNXL

MACRO TLATNX4
    CLASS CORE ;
    FOREIGN TLATNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.400 1.380 10.420 3.220 ;
        RECT  10.060 1.380 10.400 3.240 ;
        RECT  10.040 1.380 10.060 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.420 9.120 1.845 ;
        RECT  9.100 2.900 9.120 3.240 ;
        RECT  8.780 1.420 9.100 3.240 ;
        RECT  8.720 1.820 8.780 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.090 0.530 2.660 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.965 1.520 5.020 1.860 ;
        RECT  4.965 2.635 5.020 2.905 ;
        RECT  4.735 1.520 4.965 2.905 ;
        RECT  4.680 1.520 4.735 1.860 ;
        RECT  4.670 2.335 4.735 2.905 ;
        RECT  4.175 2.335 4.670 2.660 ;
        RECT  3.010 2.335 4.175 2.565 ;
        RECT  2.670 2.280 3.010 2.620 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.220 0.400 ;
        RECT  10.700 -0.400 11.040 1.060 ;
        RECT  9.760 -0.400 10.700 0.400 ;
        RECT  9.420 -0.400 9.760 1.060 ;
        RECT  7.660 -0.400 9.420 0.400 ;
        RECT  7.320 -0.400 7.660 0.575 ;
        RECT  4.980 -0.400 7.320 0.400 ;
        RECT  4.640 -0.400 4.980 0.575 ;
        RECT  2.340 -0.400 4.640 0.400 ;
        RECT  2.000 -0.400 2.340 0.575 ;
        RECT  0.520 -0.400 2.000 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 4.640 11.220 5.440 ;
        RECT  10.700 4.090 11.040 5.440 ;
        RECT  9.760 4.640 10.700 5.440 ;
        RECT  9.420 4.090 9.760 5.440 ;
        RECT  8.480 4.640 9.420 5.440 ;
        RECT  8.140 4.090 8.480 5.440 ;
        RECT  7.060 4.640 8.140 5.440 ;
        RECT  6.720 4.465 7.060 5.440 ;
        RECT  4.780 4.640 6.720 5.440 ;
        RECT  4.440 4.090 4.780 5.440 ;
        RECT  2.220 4.640 4.440 5.440 ;
        RECT  1.880 4.090 2.220 5.440 ;
        RECT  0.520 4.640 1.880 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.650 2.270 10.880 3.805 ;
        RECT  8.490 3.575 10.650 3.805 ;
        RECT  8.260 1.830 8.490 3.805 ;
        RECT  7.740 1.830 8.260 2.060 ;
        RECT  7.760 3.520 8.260 3.805 ;
        RECT  7.680 2.320 8.020 2.730 ;
        RECT  6.850 3.520 7.760 3.860 ;
        RECT  7.400 1.190 7.740 2.060 ;
        RECT  6.895 2.320 7.680 2.550 ;
        RECT  7.125 1.720 7.400 2.060 ;
        RECT  6.665 0.940 6.895 2.550 ;
        RECT  6.510 2.780 6.850 3.860 ;
        RECT  6.300 0.940 6.665 1.170 ;
        RECT  6.215 2.320 6.665 2.550 ;
        RECT  6.205 1.520 6.435 1.870 ;
        RECT  5.960 0.825 6.300 1.170 ;
        RECT  5.985 2.320 6.215 4.375 ;
        RECT  5.635 1.640 6.205 1.870 ;
        RECT  5.245 4.145 5.985 4.375 ;
        RECT  3.320 0.830 5.960 1.170 ;
        RECT  5.405 1.640 5.635 3.380 ;
        RECT  4.270 3.150 5.405 3.380 ;
        RECT  5.015 3.630 5.245 4.375 ;
        RECT  3.500 3.630 5.015 3.860 ;
        RECT  4.040 2.925 4.270 3.380 ;
        RECT  3.750 2.925 4.040 3.155 ;
        RECT  3.400 2.795 3.750 3.155 ;
        RECT  3.390 1.520 3.730 1.860 ;
        RECT  3.160 3.630 3.500 4.020 ;
        RECT  1.675 2.925 3.400 3.155 ;
        RECT  2.535 1.575 3.390 1.805 ;
        RECT  2.305 0.805 2.535 1.805 ;
        RECT  1.080 0.805 2.305 1.035 ;
        RECT  1.675 1.265 1.780 1.605 ;
        RECT  1.445 1.265 1.675 3.245 ;
        RECT  1.440 1.265 1.445 1.605 ;
        RECT  1.335 2.870 1.445 3.245 ;
        RECT  1.080 1.960 1.215 2.300 ;
        RECT  0.850 0.805 1.080 3.950 ;
        RECT  0.740 1.320 0.850 1.660 ;
        RECT  0.740 3.610 0.850 3.950 ;
    END
END TLATNX4

MACRO TLATNX2
    CLASS CORE ;
    FOREIGN TLATNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.685 0.815 7.740 2.100 ;
        RECT  7.455 0.815 7.685 3.820 ;
        RECT  7.400 0.815 7.455 2.100 ;
        RECT  7.345 3.010 7.455 3.820 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.165 2.940 6.435 3.220 ;
        RECT  6.165 1.390 6.220 1.845 ;
        RECT  5.935 1.390 6.165 4.220 ;
        RECT  5.880 1.390 5.935 1.730 ;
        RECT  5.770 3.880 5.935 4.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 1.845 0.540 2.390 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 1.860 2.735 2.200 ;
        RECT  2.395 1.860 2.625 2.635 ;
        RECT  2.195 2.405 2.395 2.635 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.980 -0.400 7.920 0.400 ;
        RECT  6.640 -0.400 6.980 0.575 ;
        RECT  4.865 -0.400 6.640 0.400 ;
        RECT  4.525 -0.400 4.865 0.575 ;
        RECT  2.385 -0.400 4.525 0.400 ;
        RECT  2.045 -0.400 2.385 0.575 ;
        RECT  0.520 -0.400 2.045 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.925 4.640 7.920 5.440 ;
        RECT  6.585 4.465 6.925 5.440 ;
        RECT  5.035 4.640 6.585 5.440 ;
        RECT  4.695 4.465 5.035 5.440 ;
        RECT  2.235 4.640 4.695 5.440 ;
        RECT  1.895 3.500 2.235 5.440 ;
        RECT  0.520 4.640 1.895 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.060 2.100 7.170 2.440 ;
        RECT  6.830 0.930 7.060 2.440 ;
        RECT  5.625 0.930 6.830 1.160 ;
        RECT  5.595 0.640 5.625 1.160 ;
        RECT  5.365 0.640 5.595 3.280 ;
        RECT  5.285 0.640 5.365 0.980 ;
        RECT  4.985 1.615 5.365 1.970 ;
        RECT  5.255 2.940 5.365 3.280 ;
        RECT  4.755 2.340 5.130 2.680 ;
        RECT  4.525 0.940 4.755 4.165 ;
        RECT  3.705 0.940 4.525 1.170 ;
        RECT  3.515 3.935 4.525 4.165 ;
        RECT  4.065 1.970 4.295 3.705 ;
        RECT  3.465 1.970 4.065 2.200 ;
        RECT  3.615 3.475 4.065 3.705 ;
        RECT  3.605 2.530 3.835 3.120 ;
        RECT  3.365 0.830 3.705 1.170 ;
        RECT  1.675 2.890 3.605 3.120 ;
        RECT  3.175 3.935 3.515 4.310 ;
        RECT  3.295 1.860 3.465 2.200 ;
        RECT  3.065 1.400 3.295 2.200 ;
        RECT  2.555 1.400 3.065 1.630 ;
        RECT  2.325 0.845 2.555 1.630 ;
        RECT  1.080 0.845 2.325 1.075 ;
        RECT  1.675 1.330 1.785 1.670 ;
        RECT  1.660 1.330 1.675 3.120 ;
        RECT  1.445 1.330 1.660 4.030 ;
        RECT  1.430 2.890 1.445 4.030 ;
        RECT  1.135 3.690 1.430 4.030 ;
        RECT  1.080 1.860 1.215 2.200 ;
        RECT  0.850 0.845 1.080 3.120 ;
        RECT  0.740 1.240 0.850 1.580 ;
        RECT  0.740 2.780 0.850 3.120 ;
    END
END TLATNX2

MACRO TLATNX1
    CLASS CORE ;
    FOREIGN TLATNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.040 1.255 7.045 3.245 ;
        RECT  6.815 1.200 7.040 3.300 ;
        RECT  6.700 1.200 6.815 1.540 ;
        RECT  6.700 2.960 6.815 3.300 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.155 0.865 6.385 3.755 ;
        RECT  6.080 0.865 6.155 1.285 ;
        RECT  5.580 3.525 6.155 3.755 ;
        RECT  5.745 0.865 6.080 1.095 ;
        RECT  5.520 0.765 5.745 1.095 ;
        RECT  5.350 3.525 5.580 4.140 ;
        RECT  5.515 0.710 5.520 1.095 ;
        RECT  5.180 0.710 5.515 1.050 ;
        RECT  5.240 3.800 5.350 4.140 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 1.845 0.530 2.380 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.360 2.500 2.935 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.400 -0.400 7.260 0.400 ;
        RECT  6.060 -0.400 6.400 0.575 ;
        RECT  4.700 -0.400 6.060 0.400 ;
        RECT  4.360 -0.400 4.700 0.575 ;
        RECT  2.170 -0.400 4.360 0.400 ;
        RECT  1.830 -0.400 2.170 0.575 ;
        RECT  0.520 -0.400 1.830 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.410 4.640 7.260 5.440 ;
        RECT  6.005 4.465 6.410 5.440 ;
        RECT  4.760 4.640 6.005 5.440 ;
        RECT  4.420 4.465 4.760 5.440 ;
        RECT  2.180 4.640 4.420 5.440 ;
        RECT  1.840 3.720 2.180 5.440 ;
        RECT  0.520 4.640 1.840 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.670 2.100 5.780 2.440 ;
        RECT  5.580 1.545 5.670 3.175 ;
        RECT  5.440 1.490 5.580 3.175 ;
        RECT  5.240 1.490 5.440 1.830 ;
        RECT  5.240 2.810 5.440 3.175 ;
        RECT  4.815 2.945 5.240 3.175 ;
        RECT  4.295 2.070 5.060 2.410 ;
        RECT  4.585 2.945 4.815 3.920 ;
        RECT  4.410 3.690 4.585 3.920 ;
        RECT  4.070 3.690 4.410 4.030 ;
        RECT  4.065 0.910 4.295 3.455 ;
        RECT  3.520 0.910 4.065 1.140 ;
        RECT  3.460 3.225 4.065 3.455 ;
        RECT  3.460 1.470 3.800 1.810 ;
        RECT  3.180 0.800 3.520 1.140 ;
        RECT  3.095 1.525 3.460 1.755 ;
        RECT  3.225 3.225 3.460 3.790 ;
        RECT  3.120 3.450 3.225 3.790 ;
        RECT  3.095 2.570 3.150 2.910 ;
        RECT  2.865 1.525 3.095 2.910 ;
        RECT  1.805 1.525 2.865 1.755 ;
        RECT  2.810 2.570 2.865 2.910 ;
        RECT  1.575 0.875 1.805 3.155 ;
        RECT  1.290 0.875 1.575 1.105 ;
        RECT  1.485 2.925 1.575 3.155 ;
        RECT  1.255 2.925 1.485 4.040 ;
        RECT  0.950 0.735 1.290 1.105 ;
        RECT  1.120 3.700 1.255 4.040 ;
        RECT  0.990 2.245 1.215 2.635 ;
        RECT  0.990 1.440 1.120 1.780 ;
        RECT  0.990 2.910 1.025 3.275 ;
        RECT  0.760 1.440 0.990 3.275 ;
    END
END TLATNX1

MACRO TLATXL
    CLASS CORE ;
    FOREIGN TLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 3.090 7.080 3.430 ;
        RECT  7.045 1.160 7.060 1.500 ;
        RECT  6.815 1.160 7.045 3.430 ;
        RECT  6.720 1.160 6.815 1.500 ;
        RECT  6.740 3.090 6.815 3.430 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.225 0.865 6.455 3.755 ;
        RECT  6.080 0.865 6.225 1.285 ;
        RECT  5.620 3.525 6.225 3.755 ;
        RECT  5.530 0.865 6.080 1.095 ;
        RECT  5.280 3.525 5.620 4.150 ;
        RECT  5.175 0.685 5.530 1.095 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.530 2.350 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 2.260 2.535 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.350 -0.400 7.260 0.400 ;
        RECT  6.010 -0.400 6.350 0.575 ;
        RECT  4.700 -0.400 6.010 0.400 ;
        RECT  4.360 -0.400 4.700 0.575 ;
        RECT  2.020 -0.400 4.360 0.400 ;
        RECT  1.680 -0.400 2.020 0.575 ;
        RECT  0.520 -0.400 1.680 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 4.640 7.260 5.440 ;
        RECT  5.980 4.465 6.320 5.440 ;
        RECT  4.860 4.640 5.980 5.440 ;
        RECT  4.520 4.465 4.860 5.440 ;
        RECT  2.095 4.640 4.520 5.440 ;
        RECT  1.755 3.460 2.095 5.440 ;
        RECT  0.520 4.640 1.755 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.755 2.100 5.810 2.440 ;
        RECT  5.620 1.400 5.755 3.135 ;
        RECT  5.525 1.400 5.620 3.190 ;
        RECT  5.190 1.400 5.525 1.740 ;
        RECT  5.470 2.100 5.525 2.440 ;
        RECT  5.280 2.850 5.525 3.190 ;
        RECT  4.990 2.960 5.280 3.190 ;
        RECT  4.800 2.070 5.140 2.410 ;
        RECT  4.760 2.960 4.990 3.905 ;
        RECT  4.185 2.070 4.800 2.300 ;
        RECT  4.325 3.675 4.760 3.905 ;
        RECT  3.985 3.620 4.325 3.960 ;
        RECT  4.125 2.070 4.185 3.285 ;
        RECT  3.955 0.790 4.125 3.285 ;
        RECT  3.895 0.790 3.955 2.300 ;
        RECT  3.375 3.055 3.955 3.285 ;
        RECT  3.340 0.790 3.895 1.020 ;
        RECT  3.295 2.480 3.600 2.820 ;
        RECT  3.140 3.055 3.375 3.590 ;
        RECT  3.000 0.680 3.340 1.020 ;
        RECT  3.260 1.390 3.295 2.820 ;
        RECT  3.065 1.390 3.260 2.765 ;
        RECT  3.035 3.250 3.140 3.590 ;
        RECT  2.970 1.390 3.065 1.620 ;
        RECT  2.630 1.280 2.970 1.620 ;
        RECT  1.675 1.390 2.630 1.620 ;
        RECT  1.525 0.865 1.675 3.135 ;
        RECT  1.445 0.865 1.525 3.700 ;
        RECT  1.220 0.865 1.445 1.095 ;
        RECT  1.295 2.905 1.445 3.700 ;
        RECT  1.260 3.470 1.295 3.700 ;
        RECT  0.920 3.470 1.260 3.810 ;
        RECT  0.880 0.805 1.220 1.095 ;
        RECT  1.065 2.060 1.215 2.405 ;
        RECT  1.065 1.450 1.120 1.790 ;
        RECT  0.835 1.450 1.065 3.110 ;
        RECT  0.780 1.450 0.835 1.790 ;
    END
END TLATXL

MACRO TLATX4
    CLASS CORE ;
    FOREIGN TLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.400 1.380 10.420 3.220 ;
        RECT  10.060 1.380 10.400 3.240 ;
        RECT  10.040 1.380 10.060 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.420 9.120 1.850 ;
        RECT  9.100 2.900 9.120 3.240 ;
        RECT  8.780 1.420 9.100 3.240 ;
        RECT  8.720 1.820 8.780 3.220 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.020 0.530 2.640 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.965 1.520 5.020 1.860 ;
        RECT  4.965 2.630 5.020 2.905 ;
        RECT  4.735 1.520 4.965 2.905 ;
        RECT  4.680 1.520 4.735 1.860 ;
        RECT  4.670 2.335 4.735 2.905 ;
        RECT  4.175 2.335 4.670 2.660 ;
        RECT  3.010 2.335 4.175 2.565 ;
        RECT  2.670 2.280 3.010 2.620 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.220 0.400 ;
        RECT  10.700 -0.400 11.040 1.060 ;
        RECT  9.760 -0.400 10.700 0.400 ;
        RECT  9.420 -0.400 9.760 1.060 ;
        RECT  7.660 -0.400 9.420 0.400 ;
        RECT  7.320 -0.400 7.660 0.575 ;
        RECT  4.980 -0.400 7.320 0.400 ;
        RECT  4.640 -0.400 4.980 0.575 ;
        RECT  2.340 -0.400 4.640 0.400 ;
        RECT  2.000 -0.400 2.340 0.575 ;
        RECT  0.520 -0.400 2.000 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 4.640 11.220 5.440 ;
        RECT  10.700 4.090 11.040 5.440 ;
        RECT  9.760 4.640 10.700 5.440 ;
        RECT  9.420 4.090 9.760 5.440 ;
        RECT  8.480 4.640 9.420 5.440 ;
        RECT  8.140 4.090 8.480 5.440 ;
        RECT  7.060 4.640 8.140 5.440 ;
        RECT  6.720 4.465 7.060 5.440 ;
        RECT  4.780 4.640 6.720 5.440 ;
        RECT  4.440 4.090 4.780 5.440 ;
        RECT  2.220 4.640 4.440 5.440 ;
        RECT  1.880 4.090 2.220 5.440 ;
        RECT  0.520 4.640 1.880 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.935 2.270 10.990 2.610 ;
        RECT  10.705 2.270 10.935 3.805 ;
        RECT  10.650 2.270 10.705 2.610 ;
        RECT  8.490 3.575 10.705 3.805 ;
        RECT  8.260 1.830 8.490 3.805 ;
        RECT  7.740 1.830 8.260 2.060 ;
        RECT  7.760 3.520 8.260 3.805 ;
        RECT  7.680 2.320 8.020 2.675 ;
        RECT  7.420 3.520 7.760 3.860 ;
        RECT  7.400 1.190 7.740 2.060 ;
        RECT  6.895 2.320 7.680 2.550 ;
        RECT  6.850 3.520 7.420 3.750 ;
        RECT  7.125 1.720 7.400 2.060 ;
        RECT  6.665 0.885 6.895 2.550 ;
        RECT  6.620 2.780 6.850 3.750 ;
        RECT  6.300 0.885 6.665 1.115 ;
        RECT  6.215 2.320 6.665 2.550 ;
        RECT  6.510 2.780 6.620 3.120 ;
        RECT  6.205 1.520 6.435 1.870 ;
        RECT  5.960 0.820 6.300 1.160 ;
        RECT  5.985 2.320 6.215 4.375 ;
        RECT  5.635 1.640 6.205 1.870 ;
        RECT  5.245 4.145 5.985 4.375 ;
        RECT  3.660 0.885 5.960 1.115 ;
        RECT  5.405 1.640 5.635 3.380 ;
        RECT  4.270 3.150 5.405 3.380 ;
        RECT  5.015 3.630 5.245 4.375 ;
        RECT  3.500 3.630 5.015 3.860 ;
        RECT  4.040 2.935 4.270 3.380 ;
        RECT  3.750 2.935 4.040 3.165 ;
        RECT  3.400 2.795 3.750 3.165 ;
        RECT  3.390 1.520 3.730 1.860 ;
        RECT  3.320 0.830 3.660 1.170 ;
        RECT  3.160 3.445 3.500 4.255 ;
        RECT  2.835 2.935 3.400 3.165 ;
        RECT  1.780 1.575 3.390 1.805 ;
        RECT  2.605 2.935 2.835 3.765 ;
        RECT  1.025 3.535 2.605 3.765 ;
        RECT  1.675 1.140 1.780 1.805 ;
        RECT  1.445 1.140 1.675 3.245 ;
        RECT  1.440 1.140 1.445 1.480 ;
        RECT  1.335 2.870 1.445 3.245 ;
        RECT  1.025 1.960 1.215 2.300 ;
        RECT  1.025 1.320 1.080 1.660 ;
        RECT  0.795 1.320 1.025 3.950 ;
        RECT  0.740 1.320 0.795 1.660 ;
    END
END TLATX4

MACRO TLATX2
    CLASS CORE ;
    FOREIGN TLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.475 1.200 7.705 3.300 ;
        RECT  7.345 1.200 7.475 1.540 ;
        RECT  7.345 2.960 7.475 3.300 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.055 2.940 6.435 3.220 ;
        RECT  6.055 3.880 6.110 4.220 ;
        RECT  5.825 1.390 6.055 4.220 ;
        RECT  5.770 3.880 5.825 4.220 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 1.845 0.540 2.390 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 2.160 2.735 2.500 ;
        RECT  2.395 2.160 2.680 2.695 ;
        RECT  2.195 2.405 2.395 2.695 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.925 -0.400 7.920 0.400 ;
        RECT  6.585 -0.400 6.925 0.575 ;
        RECT  4.865 -0.400 6.585 0.400 ;
        RECT  4.525 -0.400 4.865 0.575 ;
        RECT  2.385 -0.400 4.525 0.400 ;
        RECT  2.045 -0.400 2.385 0.575 ;
        RECT  0.520 -0.400 2.045 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.925 4.640 7.920 5.440 ;
        RECT  6.585 4.465 6.925 5.440 ;
        RECT  5.035 4.640 6.585 5.440 ;
        RECT  4.695 4.465 5.035 5.440 ;
        RECT  2.435 4.640 4.695 5.440 ;
        RECT  2.095 4.080 2.435 5.440 ;
        RECT  0.520 4.640 2.095 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.055 2.100 7.165 2.440 ;
        RECT  6.825 0.865 7.055 2.440 ;
        RECT  5.625 0.865 6.825 1.095 ;
        RECT  5.595 0.695 5.625 1.095 ;
        RECT  5.365 0.695 5.595 3.280 ;
        RECT  5.285 0.695 5.365 0.925 ;
        RECT  5.005 1.615 5.365 1.845 ;
        RECT  5.255 2.940 5.365 3.280 ;
        RECT  4.545 2.340 5.130 2.680 ;
        RECT  4.775 1.615 5.005 1.970 ;
        RECT  4.315 0.955 4.545 4.165 ;
        RECT  3.705 0.955 4.315 1.185 ;
        RECT  3.715 3.935 4.315 4.165 ;
        RECT  3.570 3.475 4.085 3.705 ;
        RECT  3.800 1.415 4.030 2.960 ;
        RECT  2.555 1.415 3.800 1.645 ;
        RECT  3.375 3.935 3.715 4.255 ;
        RECT  3.365 0.845 3.705 1.185 ;
        RECT  3.340 1.915 3.570 3.705 ;
        RECT  3.065 1.915 3.340 2.145 ;
        RECT  1.675 3.475 3.340 3.705 ;
        RECT  2.325 0.845 2.555 1.645 ;
        RECT  1.080 0.845 2.325 1.075 ;
        RECT  1.675 1.340 1.785 1.680 ;
        RECT  1.445 1.340 1.675 4.030 ;
        RECT  1.335 3.690 1.445 4.030 ;
        RECT  1.025 2.060 1.215 2.405 ;
        RECT  1.025 0.845 1.080 1.580 ;
        RECT  1.025 2.780 1.080 3.120 ;
        RECT  0.850 0.845 1.025 3.120 ;
        RECT  0.795 1.240 0.850 3.120 ;
        RECT  0.740 1.240 0.795 1.580 ;
        RECT  0.740 2.780 0.795 3.120 ;
    END
END TLATX2

MACRO TLATX1
    CLASS CORE ;
    FOREIGN TLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.040 1.255 7.045 2.075 ;
        RECT  6.815 1.200 7.040 3.740 ;
        RECT  6.700 1.200 6.815 1.540 ;
        RECT  6.810 1.845 6.815 3.740 ;
        RECT  6.700 2.930 6.810 3.740 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.155 0.865 6.385 3.755 ;
        RECT  6.080 0.865 6.155 1.290 ;
        RECT  5.580 3.525 6.155 3.755 ;
        RECT  5.745 0.865 6.080 1.095 ;
        RECT  5.520 0.720 5.745 1.095 ;
        RECT  5.350 3.525 5.580 4.140 ;
        RECT  5.515 0.665 5.520 1.095 ;
        RECT  5.180 0.665 5.515 1.005 ;
        RECT  5.240 3.800 5.350 4.140 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 1.845 0.530 2.380 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.380 2.570 2.955 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.400 -0.400 7.260 0.400 ;
        RECT  6.060 -0.400 6.400 0.575 ;
        RECT  4.700 -0.400 6.060 0.400 ;
        RECT  4.360 -0.400 4.700 0.575 ;
        RECT  2.170 -0.400 4.360 0.400 ;
        RECT  1.830 -0.400 2.170 0.575 ;
        RECT  0.520 -0.400 1.830 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.370 4.640 7.260 5.440 ;
        RECT  6.030 4.465 6.370 5.440 ;
        RECT  4.760 4.640 6.030 5.440 ;
        RECT  4.420 4.465 4.760 5.440 ;
        RECT  2.250 4.640 4.420 5.440 ;
        RECT  1.910 3.760 2.250 5.440 ;
        RECT  0.520 4.640 1.910 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.725 2.100 5.780 2.440 ;
        RECT  5.580 1.545 5.725 3.175 ;
        RECT  5.495 1.490 5.580 3.175 ;
        RECT  5.240 1.490 5.495 1.830 ;
        RECT  5.440 2.100 5.495 2.440 ;
        RECT  5.240 2.810 5.495 3.175 ;
        RECT  4.815 2.945 5.240 3.175 ;
        RECT  4.295 2.070 5.060 2.410 ;
        RECT  4.585 2.945 4.815 3.920 ;
        RECT  4.410 3.690 4.585 3.920 ;
        RECT  4.070 3.690 4.410 4.030 ;
        RECT  4.065 2.070 4.295 3.455 ;
        RECT  3.935 2.070 4.065 2.300 ;
        RECT  3.570 3.225 4.065 3.455 ;
        RECT  3.705 0.830 3.935 2.300 ;
        RECT  3.410 2.590 3.750 2.930 ;
        RECT  3.520 0.830 3.705 1.060 ;
        RECT  3.340 3.225 3.570 4.340 ;
        RECT  3.180 0.720 3.520 1.060 ;
        RECT  3.215 2.590 3.410 2.820 ;
        RECT  3.230 4.000 3.340 4.340 ;
        RECT  2.985 1.430 3.215 2.820 ;
        RECT  2.850 1.430 2.985 1.770 ;
        RECT  1.805 1.485 2.850 1.715 ;
        RECT  1.680 0.875 1.805 1.715 ;
        RECT  1.540 0.875 1.680 3.110 ;
        RECT  1.450 0.875 1.540 4.080 ;
        RECT  1.290 0.875 1.450 1.105 ;
        RECT  1.310 2.880 1.450 4.080 ;
        RECT  1.120 3.740 1.310 4.080 ;
        RECT  0.925 0.735 1.290 1.105 ;
        RECT  0.990 2.245 1.215 2.635 ;
        RECT  0.990 1.440 1.120 1.780 ;
        RECT  0.990 2.910 1.080 3.250 ;
        RECT  0.760 1.440 0.990 3.250 ;
        RECT  0.740 2.910 0.760 3.250 ;
    END
END TLATX1

MACRO TTLATXL
    CLASS CORE ;
    FOREIGN TTLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.265 6.190 1.495 ;
        RECT  5.625 1.265 5.855 3.825 ;
        RECT  5.455 3.485 5.625 3.825 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.550 2.240 7.125 2.685 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  7.395 2.115 7.800 2.720 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.730 2.375 2.500 2.790 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.715 -0.400 8.580 0.400 ;
        RECT  7.375 -0.400 7.715 0.575 ;
        RECT  4.630 -0.400 7.375 0.400 ;
        RECT  4.290 -0.400 4.630 0.575 ;
        RECT  2.170 -0.400 4.290 0.400 ;
        RECT  0.420 -0.400 2.170 0.575 ;
        RECT  0.000 -0.400 0.420 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.215 4.640 8.580 5.440 ;
        RECT  6.875 2.960 7.215 5.440 ;
        RECT  4.445 4.640 6.875 5.440 ;
        RECT  4.215 3.540 4.445 5.440 ;
        RECT  4.015 3.540 4.215 3.770 ;
        RECT  1.390 4.640 4.215 5.440 ;
        RECT  1.050 4.465 1.390 5.440 ;
        RECT  0.000 4.640 1.050 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.265 1.215 8.320 1.555 ;
        RECT  8.210 1.215 8.265 3.245 ;
        RECT  8.035 0.805 8.210 3.245 ;
        RECT  7.980 0.805 8.035 1.555 ;
        RECT  7.595 3.015 8.035 3.245 ;
        RECT  1.595 0.805 7.980 1.035 ;
        RECT  6.650 1.270 6.915 1.500 ;
        RECT  6.420 1.270 6.650 1.955 ;
        RECT  6.320 3.015 6.495 3.245 ;
        RECT  6.320 1.725 6.420 1.955 ;
        RECT  6.090 1.725 6.320 4.350 ;
        RECT  5.150 1.265 5.390 1.495 ;
        RECT  4.920 1.265 5.150 3.825 ;
        RECT  4.735 3.485 4.920 3.825 ;
        RECT  3.710 2.125 4.690 2.540 ;
        RECT  2.285 4.085 3.985 4.315 ;
        RECT  3.480 1.265 3.710 3.770 ;
        RECT  3.005 1.265 3.480 1.495 ;
        RECT  0.815 3.540 3.480 3.770 ;
        RECT  3.050 2.885 3.245 3.290 ;
        RECT  3.015 1.835 3.050 3.290 ;
        RECT  2.820 1.835 3.015 3.115 ;
        RECT  1.420 1.835 2.820 2.065 ;
        RECT  2.055 4.000 2.285 4.315 ;
        RECT  0.350 4.000 2.055 4.230 ;
        RECT  1.230 0.805 1.595 1.105 ;
        RECT  1.310 1.350 1.420 2.065 ;
        RECT  1.080 1.350 1.310 3.165 ;
        RECT  0.740 2.935 1.080 3.165 ;
        RECT  0.585 3.410 0.815 3.770 ;
        RECT  0.350 1.380 0.620 1.720 ;
        RECT  0.120 1.380 0.350 4.230 ;
    END
END TTLATXL

MACRO TTLATX4
    CLASS CORE ;
    FOREIGN TTLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TTLATXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  12.080 1.400 12.205 1.740 ;
        RECT  11.970 1.400 12.080 3.205 ;
        RECT  11.740 1.090 11.970 3.205 ;
        RECT  10.340 1.090 11.740 1.320 ;
        RECT  11.360 2.380 11.740 3.780 ;
        RECT  10.300 2.865 11.360 3.205 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.340 1.995 13.720 2.660 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  14.000 1.820 14.380 2.465 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 1.820 4.175 2.235 ;
        RECT  3.630 1.820 3.970 2.290 ;
        RECT  3.515 1.820 3.630 2.235 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.785 -0.400 15.180 0.400 ;
        RECT  13.555 -0.400 13.785 0.950 ;
        RECT  9.270 -0.400 13.555 0.400 ;
        RECT  8.930 -0.400 9.270 0.575 ;
        RECT  7.910 -0.400 8.930 0.400 ;
        RECT  7.570 -0.400 7.910 0.575 ;
        RECT  6.530 -0.400 7.570 0.400 ;
        RECT  6.190 -0.400 6.530 0.575 ;
        RECT  4.045 -0.400 6.190 0.400 ;
        RECT  3.705 -0.400 4.045 0.575 ;
        RECT  2.180 -0.400 3.705 0.400 ;
        RECT  1.840 -0.400 2.180 0.575 ;
        RECT  0.620 -0.400 1.840 0.400 ;
        RECT  0.280 -0.400 0.620 0.575 ;
        RECT  0.000 -0.400 0.280 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.120 4.640 15.180 5.440 ;
        RECT  13.780 3.150 14.120 5.440 ;
        RECT  9.275 4.640 13.780 5.440 ;
        RECT  8.935 4.090 9.275 5.440 ;
        RECT  7.990 4.640 8.935 5.440 ;
        RECT  7.650 4.090 7.990 5.440 ;
        RECT  5.905 4.640 7.650 5.440 ;
        RECT  5.565 4.465 5.905 5.440 ;
        RECT  3.970 4.640 5.565 5.440 ;
        RECT  3.630 4.465 3.970 5.440 ;
        RECT  1.180 4.640 3.630 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.615 1.335 14.845 4.030 ;
        RECT  14.275 0.750 14.615 1.565 ;
        RECT  14.505 2.750 14.615 4.030 ;
        RECT  13.315 1.335 14.275 1.565 ;
        RECT  13.060 3.000 13.400 4.280 ;
        RECT  13.085 0.630 13.315 1.565 ;
        RECT  9.845 0.630 13.085 0.860 ;
        RECT  12.970 3.000 13.060 3.230 ;
        RECT  12.855 2.460 12.970 3.230 ;
        RECT  12.625 1.330 12.855 3.230 ;
        RECT  12.240 4.000 12.580 4.340 ;
        RECT  9.920 4.055 12.240 4.285 ;
        RECT  11.275 1.550 11.440 1.780 ;
        RECT  11.045 1.550 11.275 1.835 ;
        RECT  9.955 1.605 11.045 1.835 ;
        RECT  9.920 1.370 9.955 1.835 ;
        RECT  9.690 1.370 9.920 4.285 ;
        RECT  9.615 0.630 9.845 1.095 ;
        RECT  9.580 1.370 9.690 3.205 ;
        RECT  5.740 0.865 9.615 1.095 ;
        RECT  6.890 1.370 9.580 1.710 ;
        RECT  7.010 2.740 9.580 3.080 ;
        RECT  7.370 2.130 9.120 2.470 ;
        RECT  6.855 2.185 7.370 2.415 ;
        RECT  6.780 2.085 6.855 2.415 ;
        RECT  6.625 2.085 6.780 3.415 ;
        RECT  6.300 4.005 6.640 4.380 ;
        RECT  6.550 1.475 6.625 3.415 ;
        RECT  6.395 1.475 6.550 2.315 ;
        RECT  5.905 3.185 6.550 3.415 ;
        RECT  5.370 1.475 6.395 1.705 ;
        RECT  5.980 2.560 6.320 2.900 ;
        RECT  6.295 4.005 6.300 4.325 ;
        RECT  0.465 4.005 6.295 4.235 ;
        RECT  5.075 2.590 5.980 2.820 ;
        RECT  5.565 3.130 5.905 3.470 ;
        RECT  5.400 0.725 5.740 1.095 ;
        RECT  4.975 3.185 5.565 3.415 ;
        RECT  1.920 0.865 5.400 1.095 ;
        RECT  5.315 1.365 5.370 1.705 ;
        RECT  5.030 1.325 5.315 1.705 ;
        RECT  5.075 1.955 5.130 2.295 ;
        RECT  4.845 1.955 5.075 2.820 ;
        RECT  2.385 1.325 5.030 1.555 ;
        RECT  4.745 3.185 4.975 3.775 ;
        RECT  4.790 1.955 4.845 2.295 ;
        RECT  2.910 2.590 4.845 2.820 ;
        RECT  2.650 3.545 4.745 3.775 ;
        RECT  2.910 1.950 2.965 2.290 ;
        RECT  2.680 1.950 2.910 2.820 ;
        RECT  2.625 1.950 2.680 2.290 ;
        RECT  1.405 2.590 2.680 2.820 ;
        RECT  2.310 3.390 2.650 3.775 ;
        RECT  0.930 3.545 2.310 3.775 ;
        RECT  1.920 1.740 1.975 2.080 ;
        RECT  1.395 3.085 1.945 3.315 ;
        RECT  1.690 0.865 1.920 2.080 ;
        RECT  1.635 1.740 1.690 2.080 ;
        RECT  1.405 1.035 1.420 1.375 ;
        RECT  1.395 1.035 1.405 2.820 ;
        RECT  1.165 1.035 1.395 3.315 ;
        RECT  1.080 1.035 1.165 1.375 ;
        RECT  0.700 2.210 0.930 3.775 ;
        RECT  0.465 1.420 0.620 1.760 ;
        RECT  0.235 1.420 0.465 4.235 ;
    END
END TTLATX4

MACRO TTLATX2
    CLASS CORE ;
    FOREIGN TTLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TTLATXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  9.165 1.420 9.240 1.760 ;
        RECT  9.165 2.810 9.240 3.195 ;
        RECT  8.935 1.420 9.165 3.195 ;
        RECT  8.900 1.420 8.935 1.760 ;
        RECT  8.900 2.635 8.935 3.195 ;
        RECT  8.795 2.965 8.900 3.195 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 2.115 11.080 2.745 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 1.820 11.740 2.435 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.950 3.940 2.290 ;
        RECT  3.515 1.845 3.745 2.290 ;
        RECT  3.130 1.950 3.515 2.290 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.500 -0.400 12.540 0.400 ;
        RECT  11.160 -0.400 11.500 0.575 ;
        RECT  7.760 -0.400 11.160 0.400 ;
        RECT  7.420 -0.400 7.760 0.575 ;
        RECT  6.150 -0.400 7.420 0.400 ;
        RECT  5.810 -0.400 6.150 0.575 ;
        RECT  3.710 -0.400 5.810 0.400 ;
        RECT  3.360 -0.400 3.710 0.905 ;
        RECT  1.320 -0.400 3.360 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.500 4.640 12.540 5.440 ;
        RECT  11.160 3.015 11.500 5.440 ;
        RECT  7.800 4.640 11.160 5.440 ;
        RECT  7.460 3.460 7.800 5.440 ;
        RECT  5.600 4.640 7.460 5.440 ;
        RECT  5.260 4.465 5.600 5.440 ;
        RECT  3.710 4.640 5.260 5.440 ;
        RECT  3.360 4.145 3.710 5.440 ;
        RECT  1.280 4.640 3.360 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.210 3.160 12.220 3.500 ;
        RECT  12.100 1.310 12.210 3.500 ;
        RECT  11.990 1.250 12.100 3.500 ;
        RECT  11.980 0.810 11.990 3.500 ;
        RECT  11.760 0.810 11.980 1.590 ;
        RECT  11.880 3.160 11.980 3.500 ;
        RECT  5.500 0.810 11.760 1.040 ;
        RECT  10.435 1.440 10.740 1.780 ;
        RECT  10.435 3.230 10.740 3.570 ;
        RECT  10.435 4.010 10.490 4.350 ;
        RECT  10.400 1.440 10.435 4.350 ;
        RECT  10.205 1.550 10.400 4.350 ;
        RECT  10.150 4.010 10.205 4.350 ;
        RECT  9.905 1.420 9.960 1.760 ;
        RECT  9.905 3.415 9.960 3.755 ;
        RECT  9.675 1.420 9.905 3.755 ;
        RECT  9.620 1.420 9.675 1.760 ;
        RECT  9.620 3.415 9.675 3.755 ;
        RECT  8.520 3.525 9.620 3.755 ;
        RECT  8.415 1.420 8.520 1.760 ;
        RECT  8.415 3.415 8.520 3.755 ;
        RECT  8.185 1.420 8.415 3.755 ;
        RECT  8.180 1.420 8.185 1.760 ;
        RECT  8.180 2.980 8.185 3.755 ;
        RECT  7.000 1.420 8.180 1.650 ;
        RECT  7.025 2.980 8.180 3.210 ;
        RECT  7.145 2.060 7.955 2.400 ;
        RECT  6.540 2.060 7.145 2.345 ;
        RECT  6.795 2.980 7.025 3.740 ;
        RECT  6.660 1.310 7.000 1.650 ;
        RECT  6.310 2.060 6.540 3.430 ;
        RECT  6.120 2.060 6.310 2.290 ;
        RECT  5.600 3.200 6.310 3.430 ;
        RECT  6.080 4.000 6.190 4.340 ;
        RECT  5.890 1.315 6.120 2.290 ;
        RECT  6.075 2.570 6.080 2.915 ;
        RECT  5.850 3.685 6.080 4.340 ;
        RECT  5.840 2.520 6.075 2.915 ;
        RECT  4.990 1.315 5.890 1.545 ;
        RECT  3.115 3.685 5.850 3.915 ;
        RECT  4.660 2.520 5.840 2.750 ;
        RECT  5.260 3.090 5.600 3.430 ;
        RECT  5.400 0.685 5.500 1.040 ;
        RECT  5.270 0.630 5.400 1.040 ;
        RECT  5.060 0.630 5.270 0.970 ;
        RECT  2.490 3.145 5.260 3.375 ;
        RECT  4.220 0.740 5.060 0.970 ;
        RECT  4.650 1.260 4.990 1.600 ;
        RECT  4.620 2.005 4.660 2.750 ;
        RECT  4.280 1.950 4.620 2.750 ;
        RECT  2.745 2.520 4.280 2.750 ;
        RECT  3.990 0.740 4.220 1.365 ;
        RECT  2.285 1.135 3.990 1.365 ;
        RECT  2.885 3.685 3.115 4.410 ;
        RECT  1.765 4.180 2.885 4.410 ;
        RECT  2.515 1.860 2.745 2.750 ;
        RECT  1.900 2.410 2.515 2.640 ;
        RECT  2.425 3.145 2.490 3.775 ;
        RECT  1.815 0.675 2.425 0.905 ;
        RECT  2.260 3.145 2.425 3.945 ;
        RECT  2.055 1.135 2.285 2.175 ;
        RECT  2.075 3.545 2.260 3.945 ;
        RECT  0.810 3.545 2.075 3.775 ;
        RECT  1.615 1.945 2.055 2.175 ;
        RECT  1.540 2.410 1.900 3.245 ;
        RECT  1.385 1.315 1.825 1.660 ;
        RECT  1.585 0.675 1.815 1.040 ;
        RECT  1.535 4.005 1.765 4.410 ;
        RECT  0.925 0.810 1.585 1.040 ;
        RECT  1.385 2.410 1.540 2.640 ;
        RECT  0.520 4.005 1.535 4.235 ;
        RECT  1.155 1.315 1.385 2.640 ;
        RECT  0.810 0.810 0.925 1.460 ;
        RECT  0.695 0.810 0.810 3.775 ;
        RECT  0.580 1.230 0.695 3.775 ;
        RECT  0.350 4.005 0.520 4.375 ;
        RECT  0.350 0.630 0.465 0.980 ;
        RECT  0.235 0.630 0.350 4.375 ;
        RECT  0.120 0.750 0.235 4.375 ;
    END
END TTLATX2

MACRO TTLATX1
    CLASS CORE ;
    FOREIGN TTLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TTLATXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.850 1.365 6.135 1.705 ;
        RECT  6.000 3.770 6.110 4.110 ;
        RECT  5.850 3.550 6.000 4.110 ;
        RECT  5.795 1.365 5.850 4.110 ;
        RECT  5.715 1.420 5.795 4.110 ;
        RECT  5.620 1.420 5.715 3.780 ;
        RECT  5.495 3.515 5.620 3.755 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.080 1.950 6.460 2.660 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  7.340 2.205 7.825 2.715 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 2.335 2.500 2.750 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.715 -0.400 8.580 0.400 ;
        RECT  7.375 -0.400 7.715 0.575 ;
        RECT  4.655 -0.400 7.375 0.400 ;
        RECT  4.315 -0.400 4.655 0.575 ;
        RECT  2.170 -0.400 4.315 0.400 ;
        RECT  0.420 -0.400 2.170 0.575 ;
        RECT  0.000 -0.400 0.420 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.570 4.640 8.580 5.440 ;
        RECT  7.230 2.960 7.570 5.440 ;
        RECT  4.750 4.640 7.230 5.440 ;
        RECT  4.520 4.010 4.750 5.440 ;
        RECT  1.825 4.640 4.520 5.440 ;
        RECT  1.485 4.465 1.825 5.440 ;
        RECT  0.000 4.640 1.485 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.210 1.215 8.320 3.300 ;
        RECT  8.090 0.805 8.210 3.300 ;
        RECT  7.980 0.805 8.090 1.555 ;
        RECT  7.950 2.960 8.090 3.300 ;
        RECT  3.860 0.805 7.980 1.035 ;
        RECT  6.700 1.270 6.925 3.300 ;
        RECT  6.700 3.990 6.720 4.330 ;
        RECT  6.695 1.270 6.700 4.330 ;
        RECT  6.575 1.270 6.695 1.500 ;
        RECT  6.470 2.960 6.695 4.330 ;
        RECT  6.380 3.990 6.470 4.330 ;
        RECT  5.360 1.485 5.390 3.000 ;
        RECT  5.160 1.370 5.360 3.000 ;
        RECT  5.130 1.370 5.160 1.715 ;
        RECT  4.235 2.125 4.910 2.470 ;
        RECT  3.935 4.030 4.275 4.370 ;
        RECT  4.005 1.365 4.235 3.770 ;
        RECT  3.150 1.365 4.005 1.595 ;
        RECT  1.375 3.540 4.005 3.770 ;
        RECT  2.285 4.085 3.935 4.315 ;
        RECT  3.520 0.750 3.860 1.090 ;
        RECT  3.620 2.950 3.730 3.290 ;
        RECT  3.390 1.900 3.620 3.290 ;
        RECT  1.595 0.805 3.520 1.035 ;
        RECT  3.070 1.900 3.390 2.130 ;
        RECT  2.785 1.845 3.070 2.130 ;
        RECT  1.420 1.845 2.785 2.075 ;
        RECT  2.055 4.000 2.285 4.315 ;
        RECT  0.630 4.000 2.055 4.230 ;
        RECT  1.230 0.805 1.595 1.105 ;
        RECT  1.400 2.810 1.455 3.150 ;
        RECT  1.400 1.350 1.420 2.075 ;
        RECT  1.170 1.350 1.400 3.150 ;
        RECT  1.145 3.460 1.375 3.770 ;
        RECT  1.080 1.350 1.170 1.690 ;
        RECT  1.115 2.810 1.170 3.150 ;
        RECT  0.815 3.460 1.145 3.690 ;
        RECT  0.585 3.350 0.815 3.690 ;
        RECT  0.350 3.945 0.630 4.285 ;
        RECT  0.350 1.380 0.620 1.720 ;
        RECT  0.120 1.380 0.350 4.285 ;
    END
END TTLATX1

MACRO TIELO
    CLASS CORE ;
    FOREIGN TIELO 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 1.470 1.105 2.100 ;
        RECT  0.800 1.200 1.080 2.100 ;
        RECT  0.740 1.200 0.800 1.540 ;
        END
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.400 1.320 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 1.320 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.780 2.740 1.120 3.080 ;
        RECT  0.530 2.740 0.780 2.970 ;
        RECT  0.300 2.010 0.530 2.970 ;
        RECT  0.190 2.010 0.300 2.350 ;
    END
END TIELO

MACRO TIEHI
    CLASS CORE ;
    FOREIGN TIEHI 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 2.405 1.105 2.635 ;
        RECT  0.850 2.405 1.080 3.645 ;
        RECT  0.800 2.660 0.850 3.645 ;
        RECT  0.740 2.835 0.800 3.645 ;
        END
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.400 1.320 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 1.320 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.780 1.010 1.120 1.350 ;
        RECT  0.550 1.120 0.780 1.350 ;
        RECT  0.320 1.120 0.550 2.360 ;
        RECT  0.210 2.020 0.320 2.360 ;
    END
END TIEHI

MACRO TBUFIXL
    CLASS CORE ;
    FOREIGN TBUFIXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 1.070 2.505 3.530 ;
        RECT  2.275 1.070 2.405 4.005 ;
        RECT  2.175 1.070 2.275 1.515 ;
        RECT  2.175 3.095 2.275 4.005 ;
        RECT  2.120 1.070 2.175 1.410 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.805 1.845 2.035 2.205 ;
        RECT  1.535 1.845 1.805 2.150 ;
        RECT  0.630 1.920 1.535 2.150 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 2.405 1.430 2.875 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.140 4.640 2.640 5.440 ;
        RECT  0.800 3.845 1.140 5.440 ;
        RECT  0.000 4.640 0.800 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.890 2.535 2.045 2.875 ;
        RECT  1.660 2.535 1.890 3.415 ;
        RECT  0.520 3.185 1.660 3.415 ;
        RECT  0.380 1.335 0.520 1.675 ;
        RECT  0.380 3.065 0.520 3.415 ;
        RECT  0.150 1.335 0.380 3.415 ;
    END
END TBUFIXL

MACRO TBUFIX8
    CLASS CORE ;
    FOREIGN TBUFIX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  7.780 1.670 8.365 3.220 ;
        RECT  7.750 1.510 7.780 3.220 ;
        RECT  6.815 1.190 7.750 3.480 ;
        RECT  6.740 1.190 6.815 1.820 ;
        RECT  5.870 3.000 6.815 3.480 ;
        RECT  5.870 1.190 6.740 1.670 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.700 2.350 3.040 2.690 ;
        RECT  2.195 2.380 2.700 2.660 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.820 1.270 2.335 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.380 -0.400 8.580 0.400 ;
        RECT  8.040 -0.400 8.380 0.575 ;
        RECT  6.980 -0.400 8.040 0.400 ;
        RECT  6.640 -0.400 6.980 0.575 ;
        RECT  5.580 -0.400 6.640 0.400 ;
        RECT  5.240 -0.400 5.580 0.575 ;
        RECT  2.720 -0.400 5.240 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  1.240 -0.400 2.380 0.400 ;
        RECT  0.900 -0.400 1.240 1.380 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.380 4.640 8.580 5.440 ;
        RECT  8.040 4.465 8.380 5.440 ;
        RECT  6.980 4.640 8.040 5.440 ;
        RECT  6.640 4.465 6.980 5.440 ;
        RECT  5.600 4.640 6.640 5.440 ;
        RECT  5.260 4.465 5.600 5.440 ;
        RECT  2.720 4.640 5.260 5.440 ;
        RECT  2.380 4.465 2.720 5.440 ;
        RECT  1.200 4.640 2.380 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.170 2.370 6.510 2.715 ;
        RECT  4.785 2.485 6.170 2.715 ;
        RECT  5.250 2.005 5.840 2.235 ;
        RECT  5.020 0.865 5.250 2.235 ;
        RECT  4.310 0.865 5.020 1.095 ;
        RECT  4.785 3.755 4.800 4.235 ;
        RECT  4.555 1.325 4.785 4.235 ;
        RECT  4.460 3.755 4.555 4.235 ;
        RECT  1.960 4.005 4.460 4.235 ;
        RECT  4.080 0.865 4.310 3.525 ;
        RECT  3.740 0.750 4.080 1.105 ;
        RECT  3.740 3.295 4.080 3.525 ;
        RECT  3.510 1.680 3.850 2.020 ;
        RECT  1.960 0.875 3.740 1.105 ;
        RECT  3.320 1.680 3.510 3.775 ;
        RECT  3.280 1.465 3.320 3.775 ;
        RECT  2.980 1.465 3.280 1.910 ;
        RECT  3.165 2.940 3.280 3.775 ;
        RECT  2.940 2.940 3.165 3.280 ;
        RECT  1.730 0.875 1.960 1.525 ;
        RECT  1.730 3.130 1.960 4.235 ;
        RECT  1.730 1.995 1.865 2.335 ;
        RECT  1.620 1.185 1.730 1.525 ;
        RECT  1.500 1.995 1.730 2.835 ;
        RECT  1.620 3.130 1.730 3.940 ;
        RECT  0.520 2.605 1.500 2.835 ;
        RECT  0.380 1.100 0.520 1.440 ;
        RECT  0.380 2.605 0.520 3.845 ;
        RECT  0.180 1.100 0.380 3.845 ;
        RECT  0.150 1.100 0.180 2.835 ;
    END
END TBUFIX8

MACRO TBUFIX4
    CLASS CORE ;
    FOREIGN TBUFIX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.260 5.800 2.660 ;
        RECT  5.420 1.260 5.740 3.230 ;
        RECT  5.400 2.890 5.420 3.230 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.790 1.280 2.130 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.900 2.090 4.110 2.320 ;
        RECT  3.670 1.845 3.900 2.320 ;
        RECT  3.430 1.845 3.670 2.125 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 -0.400 6.600 0.400 ;
        RECT  6.080 -0.400 6.420 0.955 ;
        RECT  5.100 -0.400 6.080 0.400 ;
        RECT  4.290 -0.400 5.100 0.575 ;
        RECT  1.120 -0.400 4.290 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 4.640 6.600 5.440 ;
        RECT  6.080 4.465 6.420 5.440 ;
        RECT  5.060 4.640 6.080 5.440 ;
        RECT  4.720 4.465 5.060 5.440 ;
        RECT  3.600 4.640 4.720 5.440 ;
        RECT  3.260 4.465 3.600 5.440 ;
        RECT  1.320 4.640 3.260 5.440 ;
        RECT  0.980 4.465 1.320 5.440 ;
        RECT  0.000 4.640 0.980 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.335 2.300 6.390 2.640 ;
        RECT  6.105 2.300 6.335 4.120 ;
        RECT  6.050 2.300 6.105 2.640 ;
        RECT  2.810 3.890 6.105 4.120 ;
        RECT  4.925 0.815 5.155 2.220 ;
        RECT  3.200 0.815 4.925 1.045 ;
        RECT  4.360 1.560 4.570 2.805 ;
        RECT  4.340 1.560 4.360 3.380 ;
        RECT  4.180 1.560 4.340 1.790 ;
        RECT  4.020 2.575 4.340 3.380 ;
        RECT  3.440 2.575 4.020 2.805 ;
        RECT  3.155 2.460 3.440 2.805 ;
        RECT  3.145 0.815 3.200 1.275 ;
        RECT  3.100 2.460 3.155 2.800 ;
        RECT  2.860 0.705 3.145 1.275 ;
        RECT  2.110 0.705 2.860 0.935 ;
        RECT  2.570 3.290 2.810 4.120 ;
        RECT  2.340 1.635 2.570 4.120 ;
        RECT  0.520 3.890 2.340 4.120 ;
        RECT  1.880 0.705 2.110 3.380 ;
        RECT  1.580 0.705 1.880 0.935 ;
        RECT  1.680 3.040 1.880 3.380 ;
        RECT  0.520 1.290 1.650 1.520 ;
        RECT  1.130 2.460 1.470 2.800 ;
        RECT  0.520 2.515 1.130 2.745 ;
        RECT  0.380 1.025 0.520 1.520 ;
        RECT  0.380 2.515 0.520 3.330 ;
        RECT  0.180 3.815 0.520 4.120 ;
        RECT  0.150 1.025 0.380 3.330 ;
    END
END TBUFIX4

MACRO TBUFIX3
    CLASS CORE ;
    FOREIGN TBUFIX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.725 1.820 5.800 2.660 ;
        RECT  5.725 1.100 5.740 1.440 ;
        RECT  5.725 2.990 5.740 3.330 ;
        RECT  5.495 1.100 5.725 3.330 ;
        RECT  5.400 1.100 5.495 1.440 ;
        RECT  5.420 1.820 5.495 2.660 ;
        RECT  5.400 2.990 5.495 3.330 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.790 1.280 2.130 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.800 1.790 4.140 2.130 ;
        RECT  3.440 1.820 3.800 2.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 -0.400 6.600 0.400 ;
        RECT  6.080 -0.400 6.420 0.575 ;
        RECT  5.060 -0.400 6.080 0.400 ;
        RECT  4.720 -0.400 5.060 0.575 ;
        RECT  3.740 -0.400 4.720 0.400 ;
        RECT  3.400 -0.400 3.740 0.575 ;
        RECT  1.320 -0.400 3.400 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 4.640 6.600 5.440 ;
        RECT  6.080 4.465 6.420 5.440 ;
        RECT  5.060 4.640 6.080 5.440 ;
        RECT  4.720 4.465 5.060 5.440 ;
        RECT  3.740 4.640 4.720 5.440 ;
        RECT  3.400 4.465 3.740 5.440 ;
        RECT  1.390 4.640 3.400 5.440 ;
        RECT  1.050 4.465 1.390 5.440 ;
        RECT  0.000 4.640 1.050 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.335 2.460 6.390 2.800 ;
        RECT  6.105 2.460 6.335 4.120 ;
        RECT  6.050 2.460 6.105 2.800 ;
        RECT  2.980 3.890 6.105 4.120 ;
        RECT  4.925 0.805 5.155 1.970 ;
        RECT  2.600 0.805 4.925 1.035 ;
        RECT  4.370 1.310 4.600 2.745 ;
        RECT  4.020 1.310 4.370 1.540 ;
        RECT  4.360 2.515 4.370 2.745 ;
        RECT  4.020 2.515 4.360 3.330 ;
        RECT  3.440 2.515 4.020 2.745 ;
        RECT  3.100 2.460 3.440 2.800 ;
        RECT  2.680 3.650 2.980 4.120 ;
        RECT  2.450 1.710 2.680 4.120 ;
        RECT  2.490 0.780 2.600 1.120 ;
        RECT  2.260 0.780 2.490 1.335 ;
        RECT  2.315 1.710 2.450 2.050 ;
        RECT  0.520 3.890 2.450 4.120 ;
        RECT  2.085 1.105 2.260 1.335 ;
        RECT  2.085 3.040 2.220 3.380 ;
        RECT  1.855 1.105 2.085 3.380 ;
        RECT  1.365 1.180 1.595 1.520 ;
        RECT  1.130 2.460 1.470 2.800 ;
        RECT  0.520 1.290 1.365 1.520 ;
        RECT  0.520 2.515 1.130 2.745 ;
        RECT  0.380 1.025 0.520 1.520 ;
        RECT  0.380 2.515 0.520 3.330 ;
        RECT  0.180 3.815 0.520 4.120 ;
        RECT  0.150 1.025 0.380 3.330 ;
    END
END TBUFIX3

MACRO TBUFIX2
    CLASS CORE ;
    FOREIGN TBUFIX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  2.445 1.070 2.565 3.405 ;
        RECT  2.335 1.070 2.445 4.020 ;
        RECT  2.195 1.070 2.335 1.515 ;
        RECT  2.215 3.175 2.335 4.020 ;
        RECT  2.160 1.070 2.195 1.410 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 1.845 2.075 2.200 ;
        RECT  1.535 1.845 1.845 2.145 ;
        RECT  0.630 1.915 1.535 2.145 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.860 2.405 1.490 2.870 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 3.960 0.400 ;
        RECT  3.440 -0.400 3.780 1.480 ;
        RECT  1.180 -0.400 3.440 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 4.640 3.960 5.440 ;
        RECT  3.440 3.215 3.780 5.440 ;
        RECT  1.180 4.640 3.440 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.950 2.495 2.105 2.870 ;
        RECT  1.720 2.495 1.950 3.415 ;
        RECT  0.520 3.185 1.720 3.415 ;
        RECT  0.380 1.330 0.520 1.670 ;
        RECT  0.380 3.060 0.520 3.415 ;
        RECT  0.150 1.330 0.380 3.415 ;
    END
END TBUFIX2

MACRO TBUFIX20
    CLASS CORE ;
    FOREIGN TBUFIX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  14.380 1.080 15.730 1.800 ;
        RECT  14.305 3.020 15.640 3.840 ;
        RECT  14.305 1.080 14.380 1.820 ;
        RECT  12.755 1.080 14.305 3.840 ;
        RECT  12.680 1.080 12.755 1.820 ;
        RECT  9.980 3.020 12.755 3.840 ;
        RECT  12.490 1.080 12.680 1.800 ;
        RECT  9.860 1.080 12.490 1.600 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.445 1.105 3.195 ;
        RECT  0.610 2.445 0.800 2.795 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 2.205 7.045 2.635 ;
        RECT  6.520 2.205 6.815 2.435 ;
        RECT  6.180 2.095 6.520 2.435 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 -0.400 16.500 0.400 ;
        RECT  15.980 -0.400 16.320 0.575 ;
        RECT  14.960 -0.400 15.980 0.400 ;
        RECT  14.620 -0.400 14.960 0.575 ;
        RECT  13.600 -0.400 14.620 0.400 ;
        RECT  13.260 -0.400 13.600 0.575 ;
        RECT  12.240 -0.400 13.260 0.400 ;
        RECT  11.900 -0.400 12.240 0.575 ;
        RECT  10.880 -0.400 11.900 0.400 ;
        RECT  10.540 -0.400 10.880 0.575 ;
        RECT  9.520 -0.400 10.540 0.400 ;
        RECT  9.180 -0.400 9.520 0.575 ;
        RECT  8.160 -0.400 9.180 0.400 ;
        RECT  7.820 -0.400 8.160 0.575 ;
        RECT  6.800 -0.400 7.820 0.400 ;
        RECT  6.460 -0.400 6.800 0.575 ;
        RECT  5.420 -0.400 6.460 0.400 ;
        RECT  5.080 -0.400 5.420 0.575 ;
        RECT  2.720 -0.400 5.080 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  1.240 -0.400 2.380 0.400 ;
        RECT  0.900 -0.400 1.240 1.450 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 4.640 16.500 5.440 ;
        RECT  15.980 4.465 16.320 5.440 ;
        RECT  15.000 4.640 15.980 5.440 ;
        RECT  14.660 4.070 15.000 5.440 ;
        RECT  13.660 4.640 14.660 5.440 ;
        RECT  13.320 4.465 13.660 5.440 ;
        RECT  12.300 4.640 13.320 5.440 ;
        RECT  11.960 4.465 12.300 5.440 ;
        RECT  10.970 4.640 11.960 5.440 ;
        RECT  10.630 4.070 10.970 5.440 ;
        RECT  9.680 4.640 10.630 5.440 ;
        RECT  9.340 4.070 9.680 5.440 ;
        RECT  8.240 4.640 9.340 5.440 ;
        RECT  7.900 4.070 8.240 5.440 ;
        RECT  6.790 4.640 7.900 5.440 ;
        RECT  6.450 4.090 6.790 5.440 ;
        RECT  5.470 4.640 6.450 5.440 ;
        RECT  5.130 4.465 5.470 5.440 ;
        RECT  2.720 4.640 5.130 5.440 ;
        RECT  2.380 4.465 2.720 5.440 ;
        RECT  1.240 4.640 2.380 5.440 ;
        RECT  0.900 3.685 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.120 2.260 12.120 2.740 ;
        RECT  9.605 2.400 11.120 2.740 ;
        RECT  9.490 1.830 10.430 2.170 ;
        RECT  9.265 2.400 9.605 3.270 ;
        RECT  9.150 1.310 9.490 2.170 ;
        RECT  8.960 2.930 9.265 3.270 ;
        RECT  7.375 1.310 9.150 1.650 ;
        RECT  8.620 2.930 8.960 4.015 ;
        RECT  7.635 1.970 8.685 2.310 ;
        RECT  8.565 2.930 8.620 3.840 ;
        RECT  4.710 3.490 8.565 3.840 ;
        RECT  7.405 1.970 7.635 3.120 ;
        RECT  6.030 2.890 7.405 3.120 ;
        RECT  7.145 0.805 7.375 1.650 ;
        RECT  4.665 0.805 7.145 1.035 ;
        RECT  7.140 1.310 7.145 1.650 ;
        RECT  5.920 1.440 6.040 1.780 ;
        RECT  5.920 2.760 6.030 3.120 ;
        RECT  5.690 1.440 5.920 3.120 ;
        RECT  4.480 1.855 4.710 3.840 ;
        RECT  4.435 0.675 4.665 1.520 ;
        RECT  4.205 1.855 4.480 2.085 ;
        RECT  1.620 3.490 4.480 3.840 ;
        RECT  3.280 0.675 4.435 0.905 ;
        RECT  3.975 1.180 4.205 2.085 ;
        RECT  3.940 2.870 4.050 3.210 ;
        RECT  3.660 1.180 3.975 1.520 ;
        RECT  3.745 2.315 3.940 3.210 ;
        RECT  3.710 1.750 3.745 3.210 ;
        RECT  3.515 1.750 3.710 2.545 ;
        RECT  3.280 1.750 3.515 1.980 ;
        RECT  3.050 0.675 3.280 1.980 ;
        RECT  3.015 2.330 3.245 2.680 ;
        RECT  2.920 1.160 3.050 1.500 ;
        RECT  2.665 2.330 3.015 2.560 ;
        RECT  1.960 1.215 2.920 1.445 ;
        RECT  2.435 1.915 2.665 2.560 ;
        RECT  0.520 1.915 2.435 2.145 ;
        RECT  1.620 1.160 1.960 1.500 ;
        RECT  0.380 1.220 0.520 2.145 ;
        RECT  0.380 3.335 0.520 3.675 ;
        RECT  0.150 1.220 0.380 3.675 ;
    END
END TBUFIX20

MACRO TBUFIX1
    CLASS CORE ;
    FOREIGN TBUFIX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 1.070 2.505 3.530 ;
        RECT  2.275 1.070 2.405 4.000 ;
        RECT  2.175 1.070 2.275 1.515 ;
        RECT  2.175 3.150 2.275 4.000 ;
        RECT  2.120 1.070 2.175 1.410 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.805 1.840 2.035 2.185 ;
        RECT  1.765 1.840 1.805 2.130 ;
        RECT  1.535 1.845 1.765 2.130 ;
        RECT  0.630 1.900 1.535 2.130 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 2.405 1.430 2.855 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.140 4.640 2.640 5.440 ;
        RECT  0.800 3.825 1.140 5.440 ;
        RECT  0.000 4.640 0.800 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.890 2.495 2.045 2.855 ;
        RECT  1.660 2.495 1.890 3.415 ;
        RECT  0.520 3.185 1.660 3.415 ;
        RECT  0.380 1.315 0.520 1.655 ;
        RECT  0.380 3.045 0.520 3.415 ;
        RECT  0.150 1.315 0.380 3.415 ;
    END
END TBUFIX1

MACRO TBUFIX16
    CLASS CORE ;
    FOREIGN TBUFIX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  11.080 1.095 11.770 1.800 ;
        RECT  11.080 2.840 11.700 3.530 ;
        RECT  11.005 1.095 11.080 1.820 ;
        RECT  11.005 2.660 11.080 3.530 ;
        RECT  9.455 1.095 11.005 3.840 ;
        RECT  9.380 1.095 9.455 1.855 ;
        RECT  9.380 2.630 9.455 3.530 ;
        RECT  7.090 1.095 9.380 1.615 ;
        RECT  7.340 2.840 9.380 3.530 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.525 1.105 3.195 ;
        RECT  0.610 2.525 0.800 2.875 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.800 1.970 5.910 2.310 ;
        RECT  5.495 1.970 5.800 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 -0.400 12.540 0.400 ;
        RECT  12.020 -0.400 12.360 0.575 ;
        RECT  11.000 -0.400 12.020 0.400 ;
        RECT  10.660 -0.400 11.000 0.575 ;
        RECT  9.560 -0.400 10.660 0.400 ;
        RECT  9.220 -0.400 9.560 0.575 ;
        RECT  8.200 -0.400 9.220 0.400 ;
        RECT  7.860 -0.400 8.200 0.575 ;
        RECT  6.840 -0.400 7.860 0.400 ;
        RECT  6.500 -0.400 6.840 0.575 ;
        RECT  5.480 -0.400 6.500 0.400 ;
        RECT  5.140 -0.400 5.480 0.575 ;
        RECT  4.100 -0.400 5.140 0.400 ;
        RECT  3.760 -0.400 4.100 0.575 ;
        RECT  1.240 -0.400 3.760 0.400 ;
        RECT  0.900 -0.400 1.240 1.450 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 4.640 12.540 5.440 ;
        RECT  12.020 4.090 12.360 5.440 ;
        RECT  11.020 4.640 12.020 5.440 ;
        RECT  10.680 4.465 11.020 5.440 ;
        RECT  9.660 4.640 10.680 5.440 ;
        RECT  9.320 4.465 9.660 5.440 ;
        RECT  8.330 4.640 9.320 5.440 ;
        RECT  7.990 4.090 8.330 5.440 ;
        RECT  7.000 4.640 7.990 5.440 ;
        RECT  6.660 4.465 7.000 5.440 ;
        RECT  5.760 4.640 6.660 5.440 ;
        RECT  5.420 4.465 5.760 5.440 ;
        RECT  4.280 4.640 5.420 5.440 ;
        RECT  3.940 3.595 4.280 5.440 ;
        RECT  1.290 4.640 3.940 5.440 ;
        RECT  0.930 4.465 1.290 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.205 2.210 9.145 2.550 ;
        RECT  6.960 2.320 8.205 2.550 ;
        RECT  6.860 1.845 7.840 2.075 ;
        RECT  6.730 2.320 6.960 3.745 ;
        RECT  6.630 0.855 6.860 2.075 ;
        RECT  5.000 3.515 6.730 3.745 ;
        RECT  4.800 0.855 6.630 1.085 ;
        RECT  6.170 1.315 6.400 3.270 ;
        RECT  5.260 1.315 6.170 1.545 ;
        RECT  5.980 2.930 6.170 3.270 ;
        RECT  5.030 1.315 5.260 2.150 ;
        RECT  4.725 1.920 5.030 2.150 ;
        RECT  4.945 3.205 5.000 4.015 ;
        RECT  4.660 3.000 4.945 4.015 ;
        RECT  4.570 0.855 4.800 1.520 ;
        RECT  3.915 1.920 4.725 2.310 ;
        RECT  3.560 3.000 4.660 3.230 ;
        RECT  4.460 1.180 4.570 1.520 ;
        RECT  3.420 1.235 4.460 1.465 ;
        RECT  3.375 3.000 3.560 3.550 ;
        RECT  3.310 1.180 3.420 1.520 ;
        RECT  3.145 1.855 3.375 3.775 ;
        RECT  3.080 0.675 3.310 1.520 ;
        RECT  1.935 4.180 3.190 4.410 ;
        RECT  2.830 1.855 3.145 2.085 ;
        RECT  2.070 3.545 3.145 3.775 ;
        RECT  2.105 0.675 3.080 0.905 ;
        RECT  2.730 2.975 2.840 3.315 ;
        RECT  2.600 1.180 2.830 2.085 ;
        RECT  2.500 2.865 2.730 3.315 ;
        RECT  2.360 1.180 2.600 1.520 ;
        RECT  2.105 2.865 2.500 3.095 ;
        RECT  1.875 0.675 2.105 3.095 ;
        RECT  1.730 3.435 2.070 3.775 ;
        RECT  1.705 4.005 1.935 4.410 ;
        RECT  1.640 0.960 1.875 1.300 ;
        RECT  0.520 4.005 1.705 4.235 ;
        RECT  0.520 1.915 1.480 2.145 ;
        RECT  0.380 1.220 0.520 2.145 ;
        RECT  0.380 3.100 0.520 4.235 ;
        RECT  0.290 1.220 0.380 4.235 ;
        RECT  0.180 1.220 0.290 3.910 ;
        RECT  0.150 1.220 0.180 3.675 ;
    END
END TBUFIX16

MACRO TBUFIX12
    CLASS CORE ;
    FOREIGN TBUFIX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  10.490 1.615 11.005 3.780 ;
        RECT  9.455 1.095 10.490 3.780 ;
        RECT  9.380 1.095 9.455 1.820 ;
        RECT  9.380 2.660 9.455 3.500 ;
        RECT  7.090 1.095 9.380 1.615 ;
        RECT  7.300 2.840 9.380 3.360 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.280 1.130 3.220 ;
        RECT  0.680 2.280 0.795 2.750 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.800 2.170 5.900 2.510 ;
        RECT  5.495 1.820 5.800 2.510 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.220 0.400 ;
        RECT  10.700 -0.400 11.040 0.575 ;
        RECT  9.620 -0.400 10.700 0.400 ;
        RECT  9.280 -0.400 9.620 0.575 ;
        RECT  8.220 -0.400 9.280 0.400 ;
        RECT  7.880 -0.400 8.220 0.575 ;
        RECT  6.840 -0.400 7.880 0.400 ;
        RECT  6.500 -0.400 6.840 0.575 ;
        RECT  5.460 -0.400 6.500 0.400 ;
        RECT  5.120 -0.400 5.460 0.575 ;
        RECT  4.090 -0.400 5.120 0.400 ;
        RECT  3.750 -0.400 4.090 0.575 ;
        RECT  1.240 -0.400 3.750 0.400 ;
        RECT  0.900 -0.400 1.240 1.410 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 4.640 11.220 5.440 ;
        RECT  10.700 4.465 11.040 5.440 ;
        RECT  9.680 4.640 10.700 5.440 ;
        RECT  9.340 4.465 9.680 5.440 ;
        RECT  8.320 4.640 9.340 5.440 ;
        RECT  7.980 4.465 8.320 5.440 ;
        RECT  6.960 4.640 7.980 5.440 ;
        RECT  6.620 4.465 6.960 5.440 ;
        RECT  5.660 4.640 6.620 5.440 ;
        RECT  5.320 3.940 5.660 5.440 ;
        RECT  4.220 4.640 5.320 5.440 ;
        RECT  3.880 3.940 4.220 5.440 ;
        RECT  1.290 4.640 3.880 5.440 ;
        RECT  0.930 4.465 1.290 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.825 2.210 8.765 2.550 ;
        RECT  6.840 2.320 7.825 2.550 ;
        RECT  6.840 1.845 7.495 2.075 ;
        RECT  6.610 0.850 6.840 2.075 ;
        RECT  6.610 2.320 6.840 3.710 ;
        RECT  4.780 0.850 6.610 1.080 ;
        RECT  4.940 3.480 6.610 3.710 ;
        RECT  6.150 1.355 6.380 3.250 ;
        RECT  5.800 1.355 6.150 1.585 ;
        RECT  6.040 2.740 6.150 3.250 ;
        RECT  5.265 2.740 6.040 2.970 ;
        RECT  5.035 2.440 5.265 2.970 ;
        RECT  4.940 2.440 5.035 2.670 ;
        RECT  3.700 2.330 4.940 2.670 ;
        RECT  4.600 3.205 4.940 4.015 ;
        RECT  4.550 0.850 4.780 1.640 ;
        RECT  3.490 3.265 4.600 3.495 ;
        RECT  4.440 1.300 4.550 1.640 ;
        RECT  3.400 1.355 4.440 1.585 ;
        RECT  3.375 3.210 3.490 3.550 ;
        RECT  3.290 1.300 3.400 1.640 ;
        RECT  3.145 2.110 3.375 3.775 ;
        RECT  3.060 0.675 3.290 1.640 ;
        RECT  2.830 2.110 3.145 2.340 ;
        RECT  2.040 3.545 3.145 3.775 ;
        RECT  1.935 4.180 3.130 4.410 ;
        RECT  2.105 0.675 3.060 0.905 ;
        RECT  2.600 1.180 2.830 2.340 ;
        RECT  2.650 2.975 2.760 3.315 ;
        RECT  2.420 2.605 2.650 3.315 ;
        RECT  2.340 1.180 2.600 1.520 ;
        RECT  2.105 2.605 2.420 2.835 ;
        RECT  1.875 0.675 2.105 2.835 ;
        RECT  1.700 3.435 2.040 3.775 ;
        RECT  1.705 4.005 1.935 4.410 ;
        RECT  1.620 1.000 1.875 1.340 ;
        RECT  0.520 4.005 1.705 4.235 ;
        RECT  0.520 1.675 1.480 1.905 ;
        RECT  0.380 1.050 0.520 1.905 ;
        RECT  0.380 3.120 0.520 4.235 ;
        RECT  0.290 1.050 0.380 4.235 ;
        RECT  0.150 1.050 0.290 3.460 ;
    END
END TBUFIX12

MACRO TBUFXL
    CLASS CORE ;
    FOREIGN TBUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.190 4.440 1.530 ;
        RECT  4.175 1.190 4.405 3.500 ;
        RECT  4.100 1.190 4.175 1.530 ;
        RECT  4.065 3.160 4.175 3.500 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.615 1.820 1.200 2.260 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.540 3.745 3.195 ;
        RECT  3.240 2.540 3.440 2.770 ;
        RECT  2.900 2.430 3.240 2.770 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 -0.400 4.620 0.400 ;
        RECT  3.420 -0.400 3.760 0.575 ;
        RECT  1.320 -0.400 3.420 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 4.640 4.620 5.440 ;
        RECT  3.220 4.465 3.620 5.440 ;
        RECT  1.320 4.640 3.220 5.440 ;
        RECT  0.980 4.465 1.320 5.440 ;
        RECT  0.000 4.640 0.980 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.820 3.795 4.160 4.135 ;
        RECT  3.855 1.900 3.910 2.240 ;
        RECT  3.625 0.865 3.855 2.240 ;
        RECT  2.740 3.875 3.820 4.105 ;
        RECT  2.760 0.865 3.625 1.095 ;
        RECT  3.570 1.900 3.625 2.240 ;
        RECT  2.090 0.630 2.760 1.095 ;
        RECT  2.670 3.040 2.740 4.105 ;
        RECT  2.440 1.460 2.670 4.105 ;
        RECT  2.330 1.460 2.440 1.800 ;
        RECT  2.400 3.040 2.440 4.105 ;
        RECT  0.520 3.875 2.400 4.105 ;
        RECT  1.950 0.630 2.090 3.380 ;
        RECT  1.860 0.865 1.950 3.380 ;
        RECT  1.735 3.040 1.860 3.380 ;
        RECT  1.260 1.200 1.600 1.540 ;
        RECT  1.150 2.640 1.490 2.980 ;
        RECT  0.520 1.255 1.260 1.485 ;
        RECT  0.520 2.695 1.150 2.925 ;
        RECT  0.385 0.750 0.520 1.485 ;
        RECT  0.385 2.695 0.520 3.530 ;
        RECT  0.180 3.875 0.520 4.390 ;
        RECT  0.155 0.750 0.385 3.530 ;
    END
END TBUFXL

MACRO TBUFX8
    CLASS CORE ;
    FOREIGN TBUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  7.120 1.820 7.705 3.220 ;
        RECT  7.045 1.510 7.120 3.220 ;
        RECT  6.460 1.265 7.045 3.280 ;
        RECT  6.180 1.265 6.460 3.525 ;
        RECT  6.155 1.265 6.180 3.985 ;
        RECT  6.080 1.265 6.155 1.820 ;
        RECT  6.080 2.660 6.155 3.985 ;
        RECT  5.320 1.265 6.080 1.645 ;
        RECT  5.840 2.885 6.080 3.985 ;
        RECT  4.740 2.885 5.840 3.280 ;
        RECT  4.615 2.885 4.740 3.985 ;
        RECT  4.400 2.890 4.615 3.985 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.090 1.105 3.195 ;
        RECT  0.610 2.090 0.875 2.430 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.330 2.140 3.670 2.480 ;
        RECT  3.085 2.195 3.330 2.480 ;
        RECT  2.985 2.195 3.085 2.635 ;
        RECT  2.755 2.195 2.985 3.570 ;
        RECT  1.840 3.340 2.755 3.570 ;
        RECT  1.800 3.220 1.840 3.570 ;
        RECT  1.800 2.590 1.810 2.965 ;
        RECT  1.570 2.590 1.800 3.570 ;
        RECT  1.470 2.590 1.570 2.965 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.680 -0.400 7.920 0.400 ;
        RECT  7.340 -0.400 7.680 0.950 ;
        RECT  6.300 -0.400 7.340 0.400 ;
        RECT  5.960 -0.400 6.300 0.950 ;
        RECT  4.980 -0.400 5.960 0.400 ;
        RECT  4.640 -0.400 4.980 0.575 ;
        RECT  3.460 -0.400 4.640 0.400 ;
        RECT  3.120 -0.400 3.460 0.575 ;
        RECT  1.320 -0.400 3.120 0.400 ;
        RECT  0.980 -0.400 1.320 1.400 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.960 4.640 7.920 5.440 ;
        RECT  6.620 4.410 6.960 5.440 ;
        RECT  5.460 4.640 6.620 5.440 ;
        RECT  5.120 4.050 5.460 5.440 ;
        RECT  4.020 4.640 5.120 5.440 ;
        RECT  3.680 4.050 4.020 5.440 ;
        RECT  1.280 4.640 3.680 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.085 1.875 5.420 2.105 ;
        RECT  4.855 0.995 5.085 2.105 ;
        RECT  4.220 0.995 4.855 1.225 ;
        RECT  4.130 2.240 4.500 2.580 ;
        RECT  3.880 0.940 4.220 1.280 ;
        RECT  3.900 1.670 4.130 3.660 ;
        RECT  2.760 1.670 3.900 1.900 ;
        RECT  3.445 3.430 3.900 3.660 ;
        RECT  3.220 0.995 3.880 1.225 ;
        RECT  3.215 3.430 3.445 4.075 ;
        RECT  2.990 0.805 3.220 1.225 ;
        RECT  0.520 3.845 3.215 4.075 ;
        RECT  2.190 0.805 2.990 1.035 ;
        RECT  2.530 1.265 2.760 1.900 ;
        RECT  2.420 1.265 2.530 1.495 ;
        RECT  2.295 2.130 2.525 3.110 ;
        RECT  2.190 2.130 2.295 2.360 ;
        RECT  1.960 0.805 2.190 2.360 ;
        RECT  1.700 1.060 1.960 1.400 ;
        RECT  1.565 1.840 1.675 2.180 ;
        RECT  1.335 1.630 1.565 2.180 ;
        RECT  0.520 1.630 1.335 1.860 ;
        RECT  0.380 0.960 0.520 1.860 ;
        RECT  0.180 3.790 0.520 4.130 ;
        RECT  0.380 2.820 0.465 3.160 ;
        RECT  0.150 0.960 0.380 3.160 ;
    END
END TBUFX8

MACRO TBUFX4
    CLASS CORE ;
    FOREIGN TBUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.065 1.820 5.140 3.220 ;
        RECT  4.990 1.265 5.065 3.220 ;
        RECT  4.850 1.265 4.990 3.645 ;
        RECT  4.760 1.265 4.850 4.125 ;
        RECT  4.660 1.265 4.760 1.605 ;
        RECT  4.510 2.845 4.760 4.125 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.790 1.280 2.130 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.845 3.745 2.230 ;
        RECT  3.035 2.000 3.515 2.230 ;
        RECT  2.805 2.000 3.035 2.800 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 -0.400 5.940 0.400 ;
        RECT  5.420 -0.400 5.760 0.575 ;
        RECT  4.200 -0.400 5.420 0.400 ;
        RECT  3.860 -0.400 4.200 0.575 ;
        RECT  1.320 -0.400 3.860 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.610 4.640 5.940 5.440 ;
        RECT  5.270 4.465 5.610 5.440 ;
        RECT  4.085 4.640 5.270 5.440 ;
        RECT  3.275 4.465 4.085 5.440 ;
        RECT  1.390 4.640 3.275 5.440 ;
        RECT  1.050 4.465 1.390 5.440 ;
        RECT  0.000 4.640 1.050 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.650 1.920 5.760 2.260 ;
        RECT  5.420 0.805 5.650 2.260 ;
        RECT  3.240 0.805 5.420 1.035 ;
        RECT  3.650 2.460 3.760 2.800 ;
        RECT  3.420 2.460 3.650 3.520 ;
        RECT  2.810 3.290 3.420 3.520 ;
        RECT  2.900 0.630 3.240 1.035 ;
        RECT  2.120 0.630 2.900 0.860 ;
        RECT  2.570 3.290 2.810 3.630 ;
        RECT  2.570 1.430 2.740 1.770 ;
        RECT  2.340 1.430 2.570 4.105 ;
        RECT  0.520 3.875 2.340 4.105 ;
        RECT  2.110 0.630 2.120 0.970 ;
        RECT  1.880 0.630 2.110 3.380 ;
        RECT  1.780 0.630 1.880 0.970 ;
        RECT  1.750 3.040 1.880 3.380 ;
        RECT  1.365 1.220 1.595 1.560 ;
        RECT  1.130 2.460 1.470 2.800 ;
        RECT  0.520 1.330 1.365 1.560 ;
        RECT  0.520 2.515 1.130 2.745 ;
        RECT  0.380 1.025 0.520 1.560 ;
        RECT  0.380 2.515 0.520 3.330 ;
        RECT  0.180 3.820 0.520 4.160 ;
        RECT  0.150 1.025 0.380 3.330 ;
    END
END TBUFX4

MACRO TBUFX3
    CLASS CORE ;
    FOREIGN TBUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.820 4.480 2.660 ;
        RECT  4.405 1.100 4.420 1.440 ;
        RECT  4.405 2.990 4.420 3.330 ;
        RECT  4.175 1.100 4.405 3.330 ;
        RECT  4.080 1.100 4.175 1.440 ;
        RECT  4.100 1.820 4.175 2.660 ;
        RECT  4.080 2.990 4.175 3.330 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.790 1.280 2.130 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 2.380 3.820 2.660 ;
        RECT  3.460 2.380 3.520 2.690 ;
        RECT  3.120 2.350 3.460 2.690 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 -0.400 5.280 0.400 ;
        RECT  4.760 -0.400 5.100 0.575 ;
        RECT  3.740 -0.400 4.760 0.400 ;
        RECT  3.400 -0.400 3.740 0.575 ;
        RECT  1.320 -0.400 3.400 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 4.640 5.280 5.440 ;
        RECT  4.760 4.465 5.100 5.440 ;
        RECT  3.740 4.640 4.760 5.440 ;
        RECT  3.400 4.465 3.740 5.440 ;
        RECT  1.390 4.640 3.400 5.440 ;
        RECT  1.050 4.465 1.390 5.440 ;
        RECT  0.000 4.640 1.050 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.015 2.460 5.070 2.800 ;
        RECT  4.785 2.460 5.015 4.120 ;
        RECT  4.730 2.460 4.785 2.800 ;
        RECT  2.980 3.890 4.785 4.120 ;
        RECT  3.605 1.630 3.835 1.970 ;
        RECT  3.245 1.630 3.605 1.860 ;
        RECT  3.015 1.105 3.245 1.860 ;
        RECT  2.600 1.105 3.015 1.335 ;
        RECT  2.680 3.085 2.980 4.120 ;
        RECT  2.450 1.710 2.680 4.120 ;
        RECT  2.260 0.780 2.600 1.335 ;
        RECT  2.315 1.710 2.450 2.050 ;
        RECT  0.520 3.890 2.450 4.120 ;
        RECT  2.085 1.105 2.260 1.335 ;
        RECT  2.085 3.040 2.220 3.380 ;
        RECT  1.855 1.105 2.085 3.380 ;
        RECT  1.365 1.180 1.595 1.520 ;
        RECT  1.130 2.460 1.470 2.800 ;
        RECT  0.520 1.290 1.365 1.520 ;
        RECT  0.520 2.515 1.130 2.745 ;
        RECT  0.380 1.025 0.520 1.520 ;
        RECT  0.380 2.515 0.520 3.330 ;
        RECT  0.180 3.815 0.520 4.120 ;
        RECT  0.150 1.025 0.380 3.330 ;
    END
END TBUFX3

MACRO TBUFX2
    CLASS CORE ;
    FOREIGN TBUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.350 4.440 1.845 ;
        RECT  4.175 1.350 4.405 4.250 ;
        RECT  4.100 1.350 4.175 1.845 ;
        RECT  4.065 2.970 4.175 4.250 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 1.820 1.275 2.130 ;
        RECT  0.615 1.790 0.955 2.130 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.490 3.745 3.195 ;
        RECT  3.240 2.490 3.440 2.720 ;
        RECT  2.900 2.380 3.240 2.720 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 -0.400 4.620 0.400 ;
        RECT  3.420 -0.400 3.760 0.575 ;
        RECT  1.320 -0.400 3.420 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 4.640 4.620 5.440 ;
        RECT  3.250 3.610 3.590 5.440 ;
        RECT  1.280 4.640 3.250 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.640 0.865 3.870 2.220 ;
        RECT  2.120 0.865 3.640 1.095 ;
        RECT  2.670 3.210 2.740 3.550 ;
        RECT  2.630 1.460 2.670 3.550 ;
        RECT  2.570 1.460 2.630 4.105 ;
        RECT  2.440 1.460 2.570 4.375 ;
        RECT  2.330 1.460 2.440 1.800 ;
        RECT  2.400 3.210 2.440 4.375 ;
        RECT  2.230 3.875 2.400 4.375 ;
        RECT  0.520 3.875 2.230 4.105 ;
        RECT  2.085 0.660 2.120 1.095 ;
        RECT  1.855 0.660 2.085 3.250 ;
        RECT  1.780 0.660 1.855 1.000 ;
        RECT  1.640 2.910 1.855 3.250 ;
        RECT  0.520 2.405 1.625 2.635 ;
        RECT  1.365 1.230 1.595 1.570 ;
        RECT  0.520 1.230 1.365 1.460 ;
        RECT  0.385 1.035 0.520 1.460 ;
        RECT  0.385 2.405 0.520 3.360 ;
        RECT  0.180 3.875 0.520 4.245 ;
        RECT  0.155 1.035 0.385 3.360 ;
    END
END TBUFX2

MACRO TBUFX20
    CLASS CORE ;
    FOREIGN TBUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 0.900 14.410 1.615 ;
        RECT  12.325 2.945 14.320 3.715 ;
        RECT  12.325 0.900 12.400 1.845 ;
        RECT  10.775 0.900 12.325 3.780 ;
        RECT  10.700 0.900 10.775 1.820 ;
        RECT  8.660 2.945 10.775 3.715 ;
        RECT  9.810 0.900 10.700 1.615 ;
        RECT  8.405 0.900 9.810 1.575 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.445 1.105 3.195 ;
        RECT  0.610 2.445 0.800 2.795 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.740 1.970 7.110 2.635 ;
        RECT  5.830 1.970 6.740 2.310 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.000 -0.400 15.180 0.400 ;
        RECT  14.660 -0.400 15.000 0.575 ;
        RECT  13.640 -0.400 14.660 0.400 ;
        RECT  13.300 -0.400 13.640 0.575 ;
        RECT  12.280 -0.400 13.300 0.400 ;
        RECT  11.940 -0.400 12.280 0.575 ;
        RECT  10.920 -0.400 11.940 0.400 ;
        RECT  10.580 -0.400 10.920 0.575 ;
        RECT  9.540 -0.400 10.580 0.400 ;
        RECT  9.200 -0.400 9.540 0.575 ;
        RECT  8.140 -0.400 9.200 0.400 ;
        RECT  7.800 -0.400 8.140 0.575 ;
        RECT  6.780 -0.400 7.800 0.400 ;
        RECT  6.440 -0.400 6.780 0.575 ;
        RECT  5.420 -0.400 6.440 0.400 ;
        RECT  5.080 -0.400 5.420 0.575 ;
        RECT  2.740 -0.400 5.080 0.400 ;
        RECT  2.400 -0.400 2.740 0.575 ;
        RECT  1.240 -0.400 2.400 0.400 ;
        RECT  0.900 -0.400 1.240 1.450 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.000 4.640 15.180 5.440 ;
        RECT  14.660 4.465 15.000 5.440 ;
        RECT  13.680 4.640 14.660 5.440 ;
        RECT  13.340 4.070 13.680 5.440 ;
        RECT  12.340 4.640 13.340 5.440 ;
        RECT  12.000 4.465 12.340 5.440 ;
        RECT  10.980 4.640 12.000 5.440 ;
        RECT  10.640 4.465 10.980 5.440 ;
        RECT  9.650 4.640 10.640 5.440 ;
        RECT  9.310 4.070 9.650 5.440 ;
        RECT  8.360 4.640 9.310 5.440 ;
        RECT  8.020 4.070 8.360 5.440 ;
        RECT  6.920 4.640 8.020 5.440 ;
        RECT  6.580 4.070 6.920 5.440 ;
        RECT  5.470 4.640 6.580 5.440 ;
        RECT  5.130 4.090 5.470 5.440 ;
        RECT  2.720 4.640 5.130 5.440 ;
        RECT  2.380 4.465 2.720 5.440 ;
        RECT  1.240 4.640 2.380 5.440 ;
        RECT  0.900 3.685 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.480 2.260 10.420 2.715 ;
        RECT  8.400 2.375 9.480 2.715 ;
        RECT  8.095 1.805 9.150 2.145 ;
        RECT  8.060 2.375 8.400 3.270 ;
        RECT  7.755 1.180 8.095 2.145 ;
        RECT  7.640 2.930 8.060 3.270 ;
        RECT  6.100 1.180 7.755 1.520 ;
        RECT  7.300 2.930 7.640 4.015 ;
        RECT  5.850 3.175 7.300 3.585 ;
        RECT  5.760 0.805 6.100 1.520 ;
        RECT  4.860 3.175 5.850 3.515 ;
        RECT  4.665 0.805 5.760 1.145 ;
        RECT  4.750 3.175 4.860 3.830 ;
        RECT  4.520 1.375 4.750 3.830 ;
        RECT  4.380 0.635 4.665 1.145 ;
        RECT  4.000 1.375 4.520 1.605 ;
        RECT  1.620 3.490 4.520 3.830 ;
        RECT  3.335 0.635 4.380 0.865 ;
        RECT  3.940 2.915 4.050 3.255 ;
        RECT  3.660 1.300 4.000 1.640 ;
        RECT  3.725 2.315 3.940 3.255 ;
        RECT  3.710 1.870 3.725 3.255 ;
        RECT  3.495 1.870 3.710 2.545 ;
        RECT  3.335 1.870 3.495 2.100 ;
        RECT  3.105 0.635 3.335 2.100 ;
        RECT  3.015 2.330 3.245 2.680 ;
        RECT  1.620 1.160 3.105 1.500 ;
        RECT  2.665 2.330 3.015 2.560 ;
        RECT  2.435 1.915 2.665 2.560 ;
        RECT  0.520 1.915 2.435 2.145 ;
        RECT  0.380 1.220 0.520 2.145 ;
        RECT  0.380 3.335 0.520 3.675 ;
        RECT  0.150 1.220 0.380 3.675 ;
    END
END TBUFX20

MACRO TBUFX1
    CLASS CORE ;
    FOREIGN TBUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.180 4.440 1.520 ;
        RECT  4.175 1.180 4.405 3.500 ;
        RECT  4.100 1.180 4.175 1.520 ;
        RECT  4.065 3.160 4.175 3.500 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.615 1.820 1.200 2.260 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.540 3.745 3.195 ;
        RECT  3.240 2.540 3.440 2.770 ;
        RECT  2.900 2.430 3.240 2.770 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 -0.400 4.620 0.400 ;
        RECT  3.420 -0.400 3.760 0.575 ;
        RECT  1.320 -0.400 3.420 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 4.640 4.620 5.440 ;
        RECT  3.250 4.465 3.590 5.440 ;
        RECT  1.280 4.640 3.250 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.820 3.875 4.160 4.260 ;
        RECT  3.625 0.865 3.855 2.240 ;
        RECT  2.725 3.875 3.820 4.105 ;
        RECT  2.120 0.865 3.625 1.095 ;
        RECT  2.670 3.260 2.725 4.105 ;
        RECT  2.440 1.460 2.670 4.105 ;
        RECT  2.330 1.460 2.440 1.800 ;
        RECT  2.385 3.260 2.440 4.105 ;
        RECT  0.520 3.875 2.385 4.105 ;
        RECT  2.065 0.630 2.120 1.095 ;
        RECT  1.835 0.630 2.065 3.600 ;
        RECT  1.780 0.630 1.835 0.970 ;
        RECT  1.640 3.260 1.835 3.600 ;
        RECT  1.265 2.640 1.605 2.980 ;
        RECT  1.260 1.200 1.600 1.540 ;
        RECT  0.520 2.695 1.265 2.925 ;
        RECT  0.520 1.255 1.260 1.485 ;
        RECT  0.385 0.750 0.520 1.485 ;
        RECT  0.385 2.695 0.520 3.530 ;
        RECT  0.180 3.875 0.520 4.390 ;
        RECT  0.155 0.750 0.385 3.530 ;
    END
END TBUFX1

MACRO TBUFX16
    CLASS CORE ;
    FOREIGN TBUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 1.095 10.450 1.850 ;
        RECT  10.345 2.930 10.380 3.270 ;
        RECT  8.795 1.095 10.345 3.780 ;
        RECT  8.720 1.095 8.795 1.820 ;
        RECT  8.720 2.660 8.795 3.610 ;
        RECT  5.850 1.095 8.720 1.615 ;
        RECT  8.590 2.840 8.720 3.610 ;
        RECT  6.020 2.840 8.590 3.360 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.525 1.105 3.195 ;
        RECT  0.610 2.525 0.800 2.875 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 1.970 4.940 2.310 ;
        RECT  4.100 1.970 4.480 2.635 ;
        RECT  3.700 1.970 4.100 2.310 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.220 0.400 ;
        RECT  10.700 -0.400 11.040 0.575 ;
        RECT  9.680 -0.400 10.700 0.400 ;
        RECT  9.340 -0.400 9.680 0.575 ;
        RECT  8.320 -0.400 9.340 0.400 ;
        RECT  7.980 -0.400 8.320 0.575 ;
        RECT  6.960 -0.400 7.980 0.400 ;
        RECT  6.620 -0.400 6.960 0.575 ;
        RECT  5.600 -0.400 6.620 0.400 ;
        RECT  5.260 -0.400 5.600 0.575 ;
        RECT  4.240 -0.400 5.260 0.400 ;
        RECT  3.900 -0.400 4.240 0.575 ;
        RECT  1.320 -0.400 3.900 0.400 ;
        RECT  0.980 -0.400 1.320 1.450 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 4.640 11.220 5.440 ;
        RECT  10.700 4.090 11.040 5.440 ;
        RECT  9.700 4.640 10.700 5.440 ;
        RECT  9.360 4.465 9.700 5.440 ;
        RECT  8.340 4.640 9.360 5.440 ;
        RECT  8.000 4.465 8.340 5.440 ;
        RECT  7.010 4.640 8.000 5.440 ;
        RECT  6.670 4.090 7.010 5.440 ;
        RECT  5.720 4.640 6.670 5.440 ;
        RECT  5.380 3.980 5.720 5.440 ;
        RECT  4.280 4.640 5.380 5.440 ;
        RECT  3.940 3.960 4.280 5.440 ;
        RECT  1.290 4.640 3.940 5.440 ;
        RECT  0.930 4.465 1.290 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.960 2.210 7.900 2.550 ;
        RECT  5.685 2.320 6.960 2.550 ;
        RECT  5.475 1.845 6.610 2.075 ;
        RECT  5.455 2.320 5.685 3.215 ;
        RECT  5.245 1.310 5.475 2.075 ;
        RECT  5.000 2.985 5.455 3.215 ;
        RECT  4.920 1.310 5.245 1.540 ;
        RECT  4.660 2.985 5.000 4.015 ;
        RECT  4.580 1.200 4.920 1.540 ;
        RECT  3.550 3.265 4.660 3.495 ;
        RECT  3.560 1.255 4.580 1.485 ;
        RECT  3.450 1.200 3.560 1.540 ;
        RECT  3.375 3.210 3.550 3.550 ;
        RECT  3.220 0.675 3.450 1.540 ;
        RECT  3.145 1.855 3.375 3.775 ;
        RECT  2.120 0.675 3.220 0.905 ;
        RECT  1.935 4.180 3.190 4.410 ;
        RECT  2.840 1.855 3.145 2.085 ;
        RECT  2.070 3.545 3.145 3.775 ;
        RECT  2.610 1.180 2.840 2.085 ;
        RECT  2.710 2.975 2.820 3.315 ;
        RECT  2.480 2.415 2.710 3.315 ;
        RECT  2.500 1.180 2.610 1.520 ;
        RECT  2.120 2.415 2.480 2.645 ;
        RECT  1.890 0.675 2.120 2.645 ;
        RECT  1.730 2.965 2.070 3.775 ;
        RECT  1.705 4.005 1.935 4.410 ;
        RECT  1.780 0.960 1.890 1.300 ;
        RECT  0.520 4.005 1.705 4.235 ;
        RECT  0.520 1.915 1.480 2.145 ;
        RECT  0.380 1.220 0.520 2.145 ;
        RECT  0.380 3.335 0.520 4.235 ;
        RECT  0.290 1.220 0.380 4.235 ;
        RECT  0.150 1.220 0.290 3.675 ;
    END
END TBUFX16

MACRO TBUFX12
    CLASS CORE ;
    FOREIGN TBUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 1.820 9.685 3.780 ;
        RECT  8.135 1.095 9.170 3.780 ;
        RECT  8.060 1.095 8.135 1.850 ;
        RECT  8.060 2.630 8.135 3.500 ;
        RECT  5.770 1.095 8.060 1.615 ;
        RECT  5.960 2.840 8.060 3.360 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.280 1.130 3.220 ;
        RECT  0.680 2.280 0.795 2.750 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.700 2.330 4.940 2.670 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.720 -0.400 9.900 0.400 ;
        RECT  9.380 -0.400 9.720 0.575 ;
        RECT  8.300 -0.400 9.380 0.400 ;
        RECT  7.960 -0.400 8.300 0.575 ;
        RECT  6.900 -0.400 7.960 0.400 ;
        RECT  6.560 -0.400 6.900 0.575 ;
        RECT  5.500 -0.400 6.560 0.400 ;
        RECT  5.160 -0.400 5.500 0.575 ;
        RECT  4.100 -0.400 5.160 0.400 ;
        RECT  3.760 -0.400 4.100 0.575 ;
        RECT  1.240 -0.400 3.760 0.400 ;
        RECT  0.900 -0.400 1.240 1.410 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.720 4.640 9.900 5.440 ;
        RECT  9.380 4.465 9.720 5.440 ;
        RECT  8.340 4.640 9.380 5.440 ;
        RECT  8.000 4.465 8.340 5.440 ;
        RECT  6.980 4.640 8.000 5.440 ;
        RECT  6.640 4.465 6.980 5.440 ;
        RECT  5.660 4.640 6.640 5.440 ;
        RECT  5.320 3.980 5.660 5.440 ;
        RECT  4.220 4.640 5.320 5.440 ;
        RECT  3.880 3.960 4.220 5.440 ;
        RECT  1.290 4.640 3.880 5.440 ;
        RECT  0.930 4.465 1.290 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.890 2.210 7.830 2.550 ;
        RECT  5.685 2.320 6.890 2.550 ;
        RECT  5.475 1.845 6.510 2.075 ;
        RECT  5.455 2.320 5.685 3.215 ;
        RECT  5.245 1.370 5.475 2.075 ;
        RECT  4.940 2.985 5.455 3.215 ;
        RECT  4.800 1.370 5.245 1.600 ;
        RECT  4.600 2.985 4.940 4.015 ;
        RECT  4.460 1.260 4.800 1.600 ;
        RECT  3.490 3.265 4.600 3.495 ;
        RECT  3.400 1.315 4.460 1.545 ;
        RECT  3.375 3.210 3.490 3.550 ;
        RECT  3.290 1.260 3.400 1.600 ;
        RECT  3.145 1.855 3.375 3.775 ;
        RECT  3.060 0.675 3.290 1.600 ;
        RECT  2.830 1.855 3.145 2.085 ;
        RECT  2.040 3.545 3.145 3.775 ;
        RECT  1.935 4.180 3.130 4.410 ;
        RECT  2.105 0.675 3.060 0.905 ;
        RECT  2.600 1.180 2.830 2.085 ;
        RECT  2.650 2.975 2.760 3.315 ;
        RECT  2.420 2.605 2.650 3.315 ;
        RECT  2.340 1.180 2.600 1.520 ;
        RECT  2.105 2.605 2.420 2.835 ;
        RECT  1.875 0.675 2.105 2.835 ;
        RECT  1.700 3.435 2.040 3.775 ;
        RECT  1.705 4.005 1.935 4.410 ;
        RECT  1.620 0.960 1.875 1.300 ;
        RECT  0.520 4.005 1.705 4.235 ;
        RECT  0.520 1.675 1.480 1.905 ;
        RECT  0.380 1.050 0.520 1.905 ;
        RECT  0.380 3.120 0.520 4.235 ;
        RECT  0.290 1.050 0.380 4.235 ;
        RECT  0.150 1.050 0.290 3.460 ;
    END
END TBUFX12

MACRO SEDFFTRXL
    CLASS CORE ;
    FOREIGN SEDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.080 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.595 0.630 3.125 1.085 ;
        RECT  2.525 0.630 2.595 0.970 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 2.160 1.840 2.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.495 1.105 2.075 ;
        RECT  0.800 1.440 0.980 2.075 ;
        RECT  0.640 1.440 0.800 1.780 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.525 2.405 23.545 2.635 ;
        RECT  23.340 2.395 23.525 3.320 ;
        RECT  23.340 1.365 23.395 1.705 ;
        RECT  23.295 1.365 23.340 3.320 ;
        RECT  23.110 1.365 23.295 2.635 ;
        RECT  23.055 1.365 23.110 1.705 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.865 1.420 24.900 3.250 ;
        RECT  24.845 1.285 24.865 3.250 ;
        RECT  24.670 1.285 24.845 3.305 ;
        RECT  24.550 1.285 24.670 1.705 ;
        RECT  24.615 2.930 24.670 3.305 ;
        RECT  24.495 1.365 24.550 1.705 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 1.820 8.455 2.310 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.845 6.125 2.200 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  12.035 1.845 12.985 2.075 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.115 -0.400 25.080 0.400 ;
        RECT  23.775 -0.400 24.115 1.705 ;
        RECT  22.265 -0.400 23.775 0.400 ;
        RECT  21.925 -0.400 22.265 0.575 ;
        RECT  19.500 -0.400 21.925 0.400 ;
        RECT  19.160 -0.400 19.500 0.880 ;
        RECT  16.670 -0.400 19.160 0.400 ;
        RECT  16.330 -0.400 16.670 1.215 ;
        RECT  13.960 -0.400 16.330 0.400 ;
        RECT  13.620 -0.400 13.960 1.470 ;
        RECT  12.560 -0.400 13.620 0.400 ;
        RECT  12.220 -0.400 12.560 0.575 ;
        RECT  8.845 -0.400 12.220 0.400 ;
        RECT  8.505 -0.400 8.845 0.870 ;
        RECT  5.925 -0.400 8.505 0.400 ;
        RECT  5.585 -0.400 5.925 0.575 ;
        RECT  2.295 -0.400 5.585 0.400 ;
        RECT  1.955 -0.400 2.295 0.890 ;
        RECT  0.610 -0.400 1.955 0.400 ;
        RECT  0.270 -0.400 0.610 0.575 ;
        RECT  0.000 -0.400 0.270 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.620 4.640 25.080 5.440 ;
        RECT  24.205 4.465 24.620 5.440 ;
        RECT  22.110 4.640 24.205 5.440 ;
        RECT  21.770 3.560 22.110 5.440 ;
        RECT  18.660 4.640 21.770 5.440 ;
        RECT  18.320 4.465 18.660 5.440 ;
        RECT  16.645 4.640 18.320 5.440 ;
        RECT  15.705 4.465 16.645 5.440 ;
        RECT  12.715 4.640 15.705 5.440 ;
        RECT  12.375 4.170 12.715 5.440 ;
        RECT  8.740 4.640 12.375 5.440 ;
        RECT  8.400 4.170 8.740 5.440 ;
        RECT  5.870 4.640 8.400 5.440 ;
        RECT  5.530 4.170 5.870 5.440 ;
        RECT  1.840 4.640 5.530 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  24.385 2.120 24.440 2.470 ;
        RECT  24.210 2.120 24.385 3.900 ;
        RECT  24.155 2.240 24.210 3.900 ;
        RECT  22.920 3.670 24.155 3.900 ;
        RECT  22.820 0.665 23.070 1.005 ;
        RECT  22.820 2.935 22.920 3.900 ;
        RECT  22.730 0.665 22.820 3.900 ;
        RECT  22.590 0.720 22.730 3.900 ;
        RECT  22.540 2.935 22.590 3.900 ;
        RECT  21.145 2.935 22.540 3.165 ;
        RECT  21.890 1.940 22.350 2.285 ;
        RECT  21.660 1.185 21.890 2.645 ;
        RECT  20.555 1.185 21.660 1.415 ;
        RECT  20.535 2.415 21.660 2.645 ;
        RECT  20.835 1.685 21.175 2.185 ;
        RECT  20.915 2.935 21.145 4.175 ;
        RECT  14.215 3.945 20.915 4.175 ;
        RECT  20.005 1.955 20.835 2.185 ;
        RECT  20.305 2.415 20.535 3.430 ;
        RECT  19.775 1.955 20.005 3.655 ;
        RECT  19.695 1.955 19.775 2.415 ;
        RECT  14.715 3.425 19.775 3.655 ;
        RECT  19.465 1.395 19.675 1.625 ;
        RECT  19.465 2.745 19.540 3.110 ;
        RECT  19.310 1.395 19.465 3.110 ;
        RECT  19.235 1.395 19.310 3.055 ;
        RECT  18.775 2.030 19.005 3.135 ;
        RECT  17.220 2.905 18.775 3.135 ;
        RECT  17.930 0.970 18.270 1.310 ;
        RECT  17.700 1.075 17.930 2.615 ;
        RECT  17.650 1.500 17.700 1.840 ;
        RECT  17.515 2.385 17.700 2.615 ;
        RECT  17.220 0.930 17.470 1.270 ;
        RECT  17.130 0.930 17.220 3.135 ;
        RECT  16.990 0.985 17.130 3.135 ;
        RECT  16.730 2.730 16.990 3.135 ;
        RECT  15.350 1.445 16.760 1.805 ;
        RECT  16.120 2.730 16.730 2.960 ;
        RECT  15.890 2.170 16.120 2.960 ;
        RECT  15.780 2.170 15.890 2.510 ;
        RECT  15.120 0.805 15.350 2.505 ;
        RECT  14.960 0.805 15.120 1.035 ;
        RECT  14.560 2.275 15.120 2.505 ;
        RECT  14.440 1.280 14.780 1.620 ;
        RECT  14.485 3.090 14.715 3.655 ;
        RECT  14.330 2.275 14.560 2.860 ;
        RECT  14.100 3.090 14.485 3.320 ;
        RECT  14.425 1.390 14.440 1.620 ;
        RECT  14.195 1.390 14.425 2.035 ;
        RECT  13.985 3.615 14.215 4.175 ;
        RECT  13.960 1.805 14.195 2.035 ;
        RECT  13.960 2.570 14.100 3.320 ;
        RECT  13.635 3.615 13.985 3.845 ;
        RECT  13.870 1.805 13.960 3.320 ;
        RECT  13.730 1.805 13.870 2.800 ;
        RECT  11.700 2.570 13.730 2.800 ;
        RECT  13.175 4.135 13.685 4.365 ;
        RECT  13.405 3.085 13.635 3.845 ;
        RECT  11.110 3.085 13.405 3.315 ;
        RECT  12.945 3.710 13.175 4.365 ;
        RECT  3.620 3.710 12.945 3.940 ;
        RECT  11.700 1.080 11.960 1.420 ;
        RECT  11.620 1.080 11.700 2.800 ;
        RECT  11.470 1.135 11.620 2.800 ;
        RECT  10.990 2.710 11.110 3.315 ;
        RECT  10.990 1.140 11.075 1.480 ;
        RECT  10.760 1.140 10.990 3.315 ;
        RECT  10.735 1.140 10.760 1.480 ;
        RECT  10.340 2.710 10.390 3.050 ;
        RECT  10.340 1.140 10.355 1.480 ;
        RECT  10.280 1.140 10.340 3.050 ;
        RECT  10.110 1.140 10.280 3.315 ;
        RECT  10.015 1.140 10.110 1.480 ;
        RECT  10.050 2.710 10.110 3.315 ;
        RECT  7.255 3.085 10.050 3.315 ;
        RECT  9.595 1.915 9.880 2.280 ;
        RECT  9.595 1.170 9.650 1.510 ;
        RECT  9.365 1.170 9.595 2.795 ;
        RECT  9.310 1.170 9.365 1.510 ;
        RECT  9.155 2.565 9.365 2.795 ;
        RECT  8.925 1.965 9.120 2.195 ;
        RECT  8.695 1.965 8.925 2.795 ;
        RECT  7.725 2.565 8.695 2.795 ;
        RECT  7.800 1.230 8.070 1.570 ;
        RECT  7.730 1.230 7.800 2.225 ;
        RECT  7.725 1.285 7.730 2.225 ;
        RECT  7.570 1.285 7.725 2.795 ;
        RECT  7.495 1.940 7.570 2.795 ;
        RECT  7.255 1.075 7.290 1.505 ;
        RECT  7.060 1.075 7.255 3.315 ;
        RECT  7.050 1.275 7.060 3.315 ;
        RECT  7.025 1.275 7.050 3.480 ;
        RECT  6.820 2.690 7.025 3.480 ;
        RECT  4.325 3.250 6.820 3.480 ;
        RECT  6.570 1.295 6.585 2.915 ;
        RECT  6.355 1.075 6.570 2.915 ;
        RECT  6.340 1.075 6.355 1.525 ;
        RECT  6.100 2.685 6.355 2.915 ;
        RECT  4.985 1.090 5.220 1.430 ;
        RECT  2.300 4.175 5.145 4.405 ;
        RECT  4.985 2.685 5.110 2.915 ;
        RECT  4.880 1.090 4.985 2.915 ;
        RECT  4.755 1.145 4.880 2.915 ;
        RECT  4.750 2.080 4.755 2.915 ;
        RECT  4.340 2.080 4.750 2.425 ;
        RECT  4.180 1.070 4.520 1.410 ;
        RECT  4.085 2.910 4.325 3.480 ;
        RECT  4.085 1.180 4.180 1.410 ;
        RECT  4.040 1.180 4.085 3.480 ;
        RECT  3.855 1.180 4.040 3.315 ;
        RECT  3.620 0.645 3.750 0.875 ;
        RECT  3.390 0.645 3.620 3.940 ;
        RECT  3.320 3.015 3.390 3.355 ;
        RECT  2.765 3.715 3.160 3.945 ;
        RECT  2.990 1.420 3.100 1.760 ;
        RECT  2.760 1.420 2.990 3.085 ;
        RECT  2.535 3.485 2.765 3.945 ;
        RECT  2.545 2.855 2.760 3.085 ;
        RECT  2.300 3.485 2.535 3.715 ;
        RECT  2.070 1.545 2.300 3.715 ;
        RECT  2.070 3.945 2.300 4.405 ;
        RECT  1.640 1.545 2.070 1.775 ;
        RECT  1.025 2.935 2.070 3.165 ;
        RECT  0.520 3.945 2.070 4.175 ;
        RECT  1.410 1.410 1.640 1.775 ;
        RECT  1.330 0.675 1.480 0.905 ;
        RECT  1.100 0.675 1.330 1.095 ;
        RECT  0.410 0.865 1.100 1.095 ;
        RECT  0.795 2.760 1.025 3.165 ;
        RECT  0.410 3.670 0.520 4.175 ;
        RECT  0.180 0.865 0.410 4.175 ;
    END
END SEDFFTRXL

MACRO SEDFFTRX4
    CLASS CORE ;
    FOREIGN SEDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFTRXL ;
    SIZE 27.720 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 0.630 3.160 1.085 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 2.160 1.840 2.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.495 1.105 2.075 ;
        RECT  0.800 1.440 0.980 2.075 ;
        RECT  0.640 1.440 0.800 1.780 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.940 1.420 24.990 1.845 ;
        RECT  24.940 2.635 24.955 3.135 ;
        RECT  24.560 1.420 24.940 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.260 1.420 26.290 1.820 ;
        RECT  25.880 1.420 26.260 3.220 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.025 1.820 8.450 2.310 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.845 6.125 2.200 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  12.355 1.845 12.985 2.075 ;
        RECT  12.015 1.790 12.355 2.130 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.930 -0.400 27.720 0.400 ;
        RECT  26.590 -0.400 26.930 1.000 ;
        RECT  25.640 -0.400 26.590 0.400 ;
        RECT  25.300 -0.400 25.640 1.005 ;
        RECT  24.320 -0.400 25.300 0.400 ;
        RECT  23.980 -0.400 24.320 1.000 ;
        RECT  22.820 -0.400 23.980 0.400 ;
        RECT  22.480 -0.400 22.820 0.575 ;
        RECT  20.225 -0.400 22.480 0.400 ;
        RECT  19.285 -0.400 20.225 0.900 ;
        RECT  16.675 -0.400 19.285 0.400 ;
        RECT  16.335 -0.400 16.675 1.215 ;
        RECT  13.965 -0.400 16.335 0.400 ;
        RECT  13.625 -0.400 13.965 1.470 ;
        RECT  12.650 -0.400 13.625 0.400 ;
        RECT  12.310 -0.400 12.650 0.575 ;
        RECT  8.845 -0.400 12.310 0.400 ;
        RECT  8.505 -0.400 8.845 1.090 ;
        RECT  5.925 -0.400 8.505 0.400 ;
        RECT  5.585 -0.400 5.925 0.575 ;
        RECT  2.295 -0.400 5.585 0.400 ;
        RECT  1.955 -0.400 2.295 0.890 ;
        RECT  0.610 -0.400 1.955 0.400 ;
        RECT  0.270 -0.400 0.610 0.575 ;
        RECT  0.000 -0.400 0.270 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.880 4.640 27.720 5.440 ;
        RECT  26.540 4.090 26.880 5.440 ;
        RECT  25.600 4.640 26.540 5.440 ;
        RECT  25.260 3.975 25.600 5.440 ;
        RECT  24.315 4.640 25.260 5.440 ;
        RECT  23.975 3.950 24.315 5.440 ;
        RECT  22.450 4.640 23.975 5.440 ;
        RECT  22.450 3.560 22.710 3.900 ;
        RECT  22.030 3.560 22.450 5.440 ;
        RECT  21.770 3.560 22.030 3.900 ;
        RECT  18.810 4.640 22.030 5.440 ;
        RECT  18.470 4.465 18.810 5.440 ;
        RECT  16.645 4.640 18.470 5.440 ;
        RECT  15.705 4.465 16.645 5.440 ;
        RECT  12.715 4.640 15.705 5.440 ;
        RECT  12.375 4.170 12.715 5.440 ;
        RECT  8.740 4.640 12.375 5.440 ;
        RECT  8.400 4.170 8.740 5.440 ;
        RECT  5.870 4.640 8.400 5.440 ;
        RECT  5.530 4.170 5.870 5.440 ;
        RECT  1.840 4.640 5.530 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  26.775 2.060 26.830 2.400 ;
        RECT  26.545 2.060 26.775 3.680 ;
        RECT  26.490 2.060 26.545 2.400 ;
        RECT  23.495 3.450 26.545 3.680 ;
        RECT  23.955 1.485 24.185 3.165 ;
        RECT  23.580 1.485 23.955 1.715 ;
        RECT  23.495 2.935 23.955 3.165 ;
        RECT  22.710 1.950 23.725 2.290 ;
        RECT  23.350 0.980 23.580 1.715 ;
        RECT  23.155 2.935 23.495 4.000 ;
        RECT  23.240 0.980 23.350 1.320 ;
        RECT  21.145 2.935 23.155 3.165 ;
        RECT  22.480 1.185 22.710 2.645 ;
        RECT  21.315 1.185 22.480 1.415 ;
        RECT  20.685 2.415 22.480 2.645 ;
        RECT  21.725 1.785 22.065 2.125 ;
        RECT  20.170 1.895 21.725 2.125 ;
        RECT  20.915 2.935 21.145 4.175 ;
        RECT  14.215 3.945 20.915 4.175 ;
        RECT  20.455 2.415 20.685 3.430 ;
        RECT  19.690 1.375 20.260 1.605 ;
        RECT  19.940 1.895 20.170 3.655 ;
        RECT  14.715 3.425 19.940 3.655 ;
        RECT  19.460 1.375 19.690 3.110 ;
        RECT  19.375 1.375 19.460 1.605 ;
        RECT  19.000 2.030 19.230 3.080 ;
        RECT  17.320 2.850 19.000 3.080 ;
        RECT  18.010 0.970 18.195 1.310 ;
        RECT  17.855 0.970 18.010 2.615 ;
        RECT  17.780 1.025 17.855 2.615 ;
        RECT  17.675 1.025 17.780 1.930 ;
        RECT  17.665 2.385 17.780 2.615 ;
        RECT  17.620 1.590 17.675 1.930 ;
        RECT  17.320 0.930 17.395 1.270 ;
        RECT  17.225 0.930 17.320 3.080 ;
        RECT  17.090 0.930 17.225 3.110 ;
        RECT  17.055 0.930 17.090 1.270 ;
        RECT  16.885 2.770 17.090 3.110 ;
        RECT  16.150 2.770 16.885 3.000 ;
        RECT  16.485 1.465 16.825 1.805 ;
        RECT  15.355 1.520 16.485 1.750 ;
        RECT  15.920 2.170 16.150 3.000 ;
        RECT  15.810 2.170 15.920 2.510 ;
        RECT  15.125 0.805 15.355 2.505 ;
        RECT  14.965 0.805 15.125 1.035 ;
        RECT  14.560 2.275 15.125 2.505 ;
        RECT  14.445 1.290 14.785 1.630 ;
        RECT  14.485 3.095 14.715 3.655 ;
        RECT  14.330 2.275 14.560 2.850 ;
        RECT  14.100 3.095 14.485 3.325 ;
        RECT  14.430 1.400 14.445 1.630 ;
        RECT  14.200 1.400 14.430 2.035 ;
        RECT  13.985 3.615 14.215 4.175 ;
        RECT  13.965 1.805 14.200 2.035 ;
        RECT  13.965 2.565 14.100 3.325 ;
        RECT  13.635 3.615 13.985 3.845 ;
        RECT  13.870 1.805 13.965 3.325 ;
        RECT  13.735 1.805 13.870 2.795 ;
        RECT  11.700 2.565 13.735 2.795 ;
        RECT  13.175 4.135 13.685 4.365 ;
        RECT  13.405 3.085 13.635 3.845 ;
        RECT  11.110 3.085 13.405 3.315 ;
        RECT  12.945 3.710 13.175 4.365 ;
        RECT  3.620 3.710 12.945 3.940 ;
        RECT  11.700 1.080 11.875 1.420 ;
        RECT  11.535 1.080 11.700 2.795 ;
        RECT  11.470 1.135 11.535 2.795 ;
        RECT  10.990 2.710 11.110 3.315 ;
        RECT  10.990 1.140 11.075 1.480 ;
        RECT  10.760 1.140 10.990 3.315 ;
        RECT  10.735 1.140 10.760 1.480 ;
        RECT  10.340 2.710 10.390 3.050 ;
        RECT  10.340 1.140 10.355 1.480 ;
        RECT  10.280 1.140 10.340 3.050 ;
        RECT  10.110 1.140 10.280 3.315 ;
        RECT  10.015 1.140 10.110 1.480 ;
        RECT  10.050 2.710 10.110 3.315 ;
        RECT  7.250 3.085 10.050 3.315 ;
        RECT  9.595 1.915 9.750 2.280 ;
        RECT  9.595 1.170 9.650 1.510 ;
        RECT  9.365 1.170 9.595 2.795 ;
        RECT  9.310 1.170 9.365 1.510 ;
        RECT  9.155 2.565 9.365 2.795 ;
        RECT  8.910 1.965 9.130 2.195 ;
        RECT  8.680 1.965 8.910 2.795 ;
        RECT  7.720 2.565 8.680 2.795 ;
        RECT  7.720 1.230 8.040 1.570 ;
        RECT  7.700 1.230 7.720 2.795 ;
        RECT  7.490 1.285 7.700 2.795 ;
        RECT  7.050 1.140 7.250 3.315 ;
        RECT  7.020 1.140 7.050 3.480 ;
        RECT  6.820 2.690 7.020 3.480 ;
        RECT  4.325 3.250 6.820 3.480 ;
        RECT  6.355 1.130 6.585 2.855 ;
        RECT  6.245 1.130 6.355 1.360 ;
        RECT  6.100 2.625 6.355 2.855 ;
        RECT  4.985 1.090 5.220 1.430 ;
        RECT  2.345 4.170 5.145 4.400 ;
        RECT  4.985 2.685 5.110 2.915 ;
        RECT  4.880 1.090 4.985 2.915 ;
        RECT  4.755 1.145 4.880 2.915 ;
        RECT  4.750 2.070 4.755 2.915 ;
        RECT  4.315 2.070 4.750 2.415 ;
        RECT  4.180 1.070 4.520 1.410 ;
        RECT  4.085 2.910 4.325 3.480 ;
        RECT  4.085 1.180 4.180 1.410 ;
        RECT  4.040 1.180 4.085 3.480 ;
        RECT  3.855 1.180 4.040 3.315 ;
        RECT  3.620 0.735 3.750 0.965 ;
        RECT  3.390 0.735 3.620 3.940 ;
        RECT  3.320 2.760 3.390 3.115 ;
        RECT  2.300 3.405 3.110 3.635 ;
        RECT  2.990 1.420 3.100 1.760 ;
        RECT  2.760 1.420 2.990 3.045 ;
        RECT  2.545 2.815 2.760 3.045 ;
        RECT  2.115 3.945 2.345 4.400 ;
        RECT  2.070 1.545 2.300 3.635 ;
        RECT  0.520 3.945 2.115 4.175 ;
        RECT  1.640 1.545 2.070 1.775 ;
        RECT  1.025 2.935 2.070 3.165 ;
        RECT  1.410 1.410 1.640 1.775 ;
        RECT  1.330 0.675 1.480 0.905 ;
        RECT  1.100 0.675 1.330 1.095 ;
        RECT  0.410 0.865 1.100 1.095 ;
        RECT  0.795 2.760 1.025 3.165 ;
        RECT  0.410 3.670 0.520 4.175 ;
        RECT  0.180 0.865 0.410 4.175 ;
    END
END SEDFFTRX4

MACRO SEDFFTRX2
    CLASS CORE ;
    FOREIGN SEDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFTRXL ;
    SIZE 26.400 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 0.630 3.160 1.085 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 2.160 1.840 2.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.495 1.105 2.075 ;
        RECT  0.800 1.440 0.980 2.075 ;
        RECT  0.640 1.440 0.800 1.780 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.745 2.405 24.865 2.635 ;
        RECT  24.730 1.455 24.785 1.845 ;
        RECT  24.730 2.405 24.745 3.095 ;
        RECT  24.500 1.455 24.730 3.095 ;
        RECT  24.445 1.455 24.500 1.795 ;
        RECT  24.405 2.755 24.500 3.095 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.100 1.285 26.185 1.515 ;
        RECT  26.025 1.285 26.100 3.040 ;
        RECT  25.870 1.285 26.025 3.095 ;
        RECT  25.725 1.455 25.870 1.795 ;
        RECT  25.685 2.755 25.870 3.095 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.025 1.820 8.450 2.310 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.845 6.125 2.200 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  12.100 1.845 12.985 2.075 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.425 -0.400 26.400 0.400 ;
        RECT  25.085 -0.400 25.425 1.145 ;
        RECT  23.165 -0.400 25.085 0.400 ;
        RECT  22.825 -0.400 23.165 0.575 ;
        RECT  20.380 -0.400 22.825 0.400 ;
        RECT  20.360 -0.400 20.380 0.560 ;
        RECT  19.420 -0.400 20.360 0.900 ;
        RECT  19.400 -0.400 19.420 0.560 ;
        RECT  16.810 -0.400 19.400 0.400 ;
        RECT  16.470 -0.400 16.810 1.215 ;
        RECT  14.100 -0.400 16.470 0.400 ;
        RECT  13.760 -0.400 14.100 1.470 ;
        RECT  12.735 -0.400 13.760 0.400 ;
        RECT  12.395 -0.400 12.735 0.575 ;
        RECT  8.845 -0.400 12.395 0.400 ;
        RECT  8.505 -0.400 8.845 1.090 ;
        RECT  5.925 -0.400 8.505 0.400 ;
        RECT  5.585 -0.400 5.925 0.575 ;
        RECT  2.295 -0.400 5.585 0.400 ;
        RECT  1.955 -0.400 2.295 0.890 ;
        RECT  0.610 -0.400 1.955 0.400 ;
        RECT  0.270 -0.400 0.610 0.575 ;
        RECT  0.000 -0.400 0.270 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.385 4.640 26.400 5.440 ;
        RECT  25.045 4.015 25.385 5.440 ;
        RECT  22.450 4.640 25.045 5.440 ;
        RECT  22.450 3.560 22.710 3.900 ;
        RECT  22.030 3.560 22.450 5.440 ;
        RECT  21.770 3.560 22.030 3.900 ;
        RECT  18.810 4.640 22.030 5.440 ;
        RECT  18.470 4.465 18.810 5.440 ;
        RECT  16.645 4.640 18.470 5.440 ;
        RECT  15.705 4.465 16.645 5.440 ;
        RECT  12.715 4.640 15.705 5.440 ;
        RECT  12.375 4.170 12.715 5.440 ;
        RECT  8.740 4.640 12.375 5.440 ;
        RECT  8.400 4.170 8.740 5.440 ;
        RECT  5.870 4.640 8.400 5.440 ;
        RECT  5.530 4.170 5.870 5.440 ;
        RECT  1.840 4.640 5.530 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  25.410 2.120 25.640 2.485 ;
        RECT  25.400 2.255 25.410 2.485 ;
        RECT  25.170 2.255 25.400 3.725 ;
        RECT  23.905 3.495 25.170 3.725 ;
        RECT  23.905 0.680 23.935 1.620 ;
        RECT  23.675 0.680 23.905 3.725 ;
        RECT  23.595 0.680 23.675 1.620 ;
        RECT  23.545 2.935 23.675 3.725 ;
        RECT  23.205 2.935 23.545 4.000 ;
        RECT  23.390 1.950 23.445 2.290 ;
        RECT  23.335 1.925 23.390 2.315 ;
        RECT  23.105 1.185 23.335 2.645 ;
        RECT  21.145 2.935 23.205 3.165 ;
        RECT  21.790 1.185 23.105 1.415 ;
        RECT  20.685 2.415 23.105 2.645 ;
        RECT  22.095 1.760 22.150 2.100 ;
        RECT  21.810 1.760 22.095 2.125 ;
        RECT  20.170 1.895 21.810 2.125 ;
        RECT  21.450 1.130 21.790 1.470 ;
        RECT  20.915 2.935 21.145 4.175 ;
        RECT  14.215 3.945 20.915 4.175 ;
        RECT  20.455 2.415 20.685 3.430 ;
        RECT  19.690 1.375 20.395 1.605 ;
        RECT  19.940 1.895 20.170 3.655 ;
        RECT  14.715 3.425 19.940 3.655 ;
        RECT  19.460 1.375 19.690 3.110 ;
        RECT  19.000 2.030 19.230 3.135 ;
        RECT  17.420 2.905 19.000 3.135 ;
        RECT  18.010 0.970 18.330 1.310 ;
        RECT  17.990 0.970 18.010 2.615 ;
        RECT  17.780 1.025 17.990 2.615 ;
        RECT  17.760 1.025 17.780 1.930 ;
        RECT  17.665 2.385 17.780 2.615 ;
        RECT  17.705 1.590 17.760 1.930 ;
        RECT  17.420 0.930 17.530 1.270 ;
        RECT  17.190 0.930 17.420 3.135 ;
        RECT  16.885 2.770 17.190 3.110 ;
        RECT  16.620 1.465 16.960 1.805 ;
        RECT  16.125 2.825 16.885 3.055 ;
        RECT  15.490 1.520 16.620 1.750 ;
        RECT  16.120 2.280 16.125 3.055 ;
        RECT  15.895 2.170 16.120 3.055 ;
        RECT  15.780 2.170 15.895 2.510 ;
        RECT  15.260 0.805 15.490 2.505 ;
        RECT  15.100 0.805 15.260 1.035 ;
        RECT  14.560 2.275 15.260 2.505 ;
        RECT  14.580 1.265 14.920 1.605 ;
        RECT  14.485 3.095 14.715 3.655 ;
        RECT  14.565 1.375 14.580 1.605 ;
        RECT  14.335 1.375 14.565 2.035 ;
        RECT  14.330 2.275 14.560 2.850 ;
        RECT  14.100 3.095 14.485 3.325 ;
        RECT  14.100 1.805 14.335 2.035 ;
        RECT  13.985 3.615 14.215 4.175 ;
        RECT  13.870 1.805 14.100 3.325 ;
        RECT  13.635 3.615 13.985 3.845 ;
        RECT  11.700 2.565 13.870 2.795 ;
        RECT  13.175 4.135 13.685 4.365 ;
        RECT  13.405 3.085 13.635 3.845 ;
        RECT  11.110 3.085 13.405 3.315 ;
        RECT  12.945 3.710 13.175 4.365 ;
        RECT  3.620 3.710 12.945 3.940 ;
        RECT  11.700 1.080 11.960 1.420 ;
        RECT  11.620 1.080 11.700 2.795 ;
        RECT  11.470 1.135 11.620 2.795 ;
        RECT  10.990 2.710 11.110 3.315 ;
        RECT  10.990 1.140 11.075 1.480 ;
        RECT  10.760 1.140 10.990 3.315 ;
        RECT  10.735 1.140 10.760 1.480 ;
        RECT  10.340 2.710 10.390 3.050 ;
        RECT  10.340 1.140 10.355 1.480 ;
        RECT  10.280 1.140 10.340 3.050 ;
        RECT  10.110 1.140 10.280 3.315 ;
        RECT  10.015 1.140 10.110 1.480 ;
        RECT  10.050 2.710 10.110 3.315 ;
        RECT  7.250 3.085 10.050 3.315 ;
        RECT  9.595 1.915 9.750 2.280 ;
        RECT  9.595 1.170 9.650 1.510 ;
        RECT  9.365 1.170 9.595 2.795 ;
        RECT  9.310 1.170 9.365 1.510 ;
        RECT  9.155 2.565 9.365 2.795 ;
        RECT  8.910 1.965 9.130 2.195 ;
        RECT  8.680 1.965 8.910 2.795 ;
        RECT  7.720 2.565 8.680 2.795 ;
        RECT  7.720 1.230 8.040 1.570 ;
        RECT  7.700 1.230 7.720 2.795 ;
        RECT  7.490 1.285 7.700 2.795 ;
        RECT  7.050 1.120 7.250 3.315 ;
        RECT  7.020 1.120 7.050 3.480 ;
        RECT  6.820 2.690 7.020 3.480 ;
        RECT  4.325 3.250 6.820 3.480 ;
        RECT  6.355 1.130 6.585 2.855 ;
        RECT  6.245 1.130 6.355 1.360 ;
        RECT  6.100 2.625 6.355 2.855 ;
        RECT  4.985 1.090 5.220 1.430 ;
        RECT  2.345 4.170 5.145 4.400 ;
        RECT  4.985 2.685 5.110 2.915 ;
        RECT  4.880 1.090 4.985 2.915 ;
        RECT  4.755 1.145 4.880 2.915 ;
        RECT  4.750 2.070 4.755 2.915 ;
        RECT  4.315 2.070 4.750 2.415 ;
        RECT  4.180 1.070 4.520 1.410 ;
        RECT  4.085 2.910 4.325 3.480 ;
        RECT  4.085 1.180 4.180 1.410 ;
        RECT  4.040 1.180 4.085 3.480 ;
        RECT  3.855 1.180 4.040 3.315 ;
        RECT  3.620 0.735 3.750 0.965 ;
        RECT  3.390 0.735 3.620 3.940 ;
        RECT  3.320 2.760 3.390 3.115 ;
        RECT  2.300 3.405 3.110 3.635 ;
        RECT  2.990 1.420 3.100 1.760 ;
        RECT  2.760 1.420 2.990 3.045 ;
        RECT  2.545 2.815 2.760 3.045 ;
        RECT  2.115 3.945 2.345 4.400 ;
        RECT  2.070 1.545 2.300 3.635 ;
        RECT  0.520 3.945 2.115 4.175 ;
        RECT  1.640 1.545 2.070 1.775 ;
        RECT  1.025 2.935 2.070 3.165 ;
        RECT  1.410 1.410 1.640 1.775 ;
        RECT  1.330 0.675 1.480 0.905 ;
        RECT  1.100 0.675 1.330 1.095 ;
        RECT  0.410 0.865 1.100 1.095 ;
        RECT  0.795 2.760 1.025 3.165 ;
        RECT  0.410 3.670 0.520 4.175 ;
        RECT  0.180 0.865 0.410 4.175 ;
    END
END SEDFFTRX2

MACRO SEDFFTRX1
    CLASS CORE ;
    FOREIGN SEDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFTRXL ;
    SIZE 25.740 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 0.630 3.160 1.085 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 2.160 1.840 2.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.495 1.105 2.075 ;
        RECT  0.800 1.440 0.980 2.075 ;
        RECT  0.640 1.440 0.800 1.780 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.180 1.345 24.235 1.845 ;
        RECT  24.180 2.405 24.205 3.200 ;
        RECT  23.950 1.345 24.180 3.200 ;
        RECT  23.900 1.345 23.950 1.845 ;
        RECT  23.900 2.660 23.950 3.200 ;
        RECT  23.895 1.345 23.900 1.685 ;
        RECT  23.870 2.845 23.900 3.200 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  25.485 1.285 25.560 3.165 ;
        RECT  25.330 1.285 25.485 3.275 ;
        RECT  25.220 1.285 25.330 1.685 ;
        RECT  25.145 2.935 25.330 3.275 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.025 1.820 8.450 2.310 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.845 6.125 2.200 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  12.245 1.845 12.985 2.075 ;
        RECT  11.905 1.790 12.245 2.130 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.800 -0.400 25.740 0.400 ;
        RECT  24.460 -0.400 24.800 0.575 ;
        RECT  22.760 -0.400 24.460 0.400 ;
        RECT  22.420 -0.400 22.760 0.575 ;
        RECT  20.155 -0.400 22.420 0.400 ;
        RECT  19.215 -0.400 20.155 0.900 ;
        RECT  16.670 -0.400 19.215 0.400 ;
        RECT  16.330 -0.400 16.670 1.215 ;
        RECT  14.000 -0.400 16.330 0.400 ;
        RECT  13.660 -0.400 14.000 1.470 ;
        RECT  12.700 -0.400 13.660 0.400 ;
        RECT  12.360 -0.400 12.700 0.575 ;
        RECT  8.845 -0.400 12.360 0.400 ;
        RECT  8.505 -0.400 8.845 1.090 ;
        RECT  5.925 -0.400 8.505 0.400 ;
        RECT  5.585 -0.400 5.925 0.575 ;
        RECT  2.295 -0.400 5.585 0.400 ;
        RECT  1.955 -0.400 2.295 0.890 ;
        RECT  0.610 -0.400 1.955 0.400 ;
        RECT  0.270 -0.400 0.610 0.575 ;
        RECT  0.000 -0.400 0.270 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.930 4.640 25.740 5.440 ;
        RECT  24.540 4.465 24.930 5.440 ;
        RECT  22.665 4.640 24.540 5.440 ;
        RECT  22.325 3.380 22.665 5.440 ;
        RECT  21.830 3.560 22.325 3.900 ;
        RECT  18.810 4.640 22.325 5.440 ;
        RECT  18.470 4.465 18.810 5.440 ;
        RECT  16.645 4.640 18.470 5.440 ;
        RECT  15.705 4.465 16.645 5.440 ;
        RECT  12.715 4.640 15.705 5.440 ;
        RECT  12.375 4.170 12.715 5.440 ;
        RECT  8.740 4.640 12.375 5.440 ;
        RECT  8.400 4.170 8.740 5.440 ;
        RECT  5.870 4.640 8.400 5.440 ;
        RECT  5.530 4.170 5.870 5.440 ;
        RECT  1.840 4.640 5.530 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  24.915 2.120 25.100 2.485 ;
        RECT  24.870 2.120 24.915 3.725 ;
        RECT  24.685 2.255 24.870 3.725 ;
        RECT  23.455 3.495 24.685 3.725 ;
        RECT  23.480 0.980 23.520 1.320 ;
        RECT  23.455 0.980 23.480 3.165 ;
        RECT  23.250 0.980 23.455 4.000 ;
        RECT  23.180 0.980 23.250 1.320 ;
        RECT  23.115 2.880 23.250 4.000 ;
        RECT  21.145 2.880 23.115 3.110 ;
        RECT  22.755 2.105 23.015 2.465 ;
        RECT  22.525 1.240 22.755 2.645 ;
        RECT  21.600 1.240 22.525 1.470 ;
        RECT  20.685 2.415 22.525 2.645 ;
        RECT  21.630 1.760 21.970 2.100 ;
        RECT  20.170 1.870 21.630 2.100 ;
        RECT  21.260 1.130 21.600 1.470 ;
        RECT  20.915 2.880 21.145 4.175 ;
        RECT  14.215 3.945 20.915 4.175 ;
        RECT  20.455 2.415 20.685 3.430 ;
        RECT  19.940 1.870 20.170 3.655 ;
        RECT  19.690 1.375 20.150 1.605 ;
        RECT  14.715 3.425 19.940 3.655 ;
        RECT  19.460 1.375 19.690 3.110 ;
        RECT  19.265 1.375 19.460 1.605 ;
        RECT  19.000 2.030 19.230 3.110 ;
        RECT  17.310 2.880 19.000 3.110 ;
        RECT  18.010 0.970 18.190 1.310 ;
        RECT  17.780 0.970 18.010 2.615 ;
        RECT  17.760 0.970 17.780 1.930 ;
        RECT  17.665 2.385 17.780 2.615 ;
        RECT  17.625 1.590 17.760 1.930 ;
        RECT  17.310 0.930 17.390 1.270 ;
        RECT  17.080 0.930 17.310 3.110 ;
        RECT  17.050 0.930 17.080 1.270 ;
        RECT  16.885 2.770 17.080 3.110 ;
        RECT  16.125 2.770 16.885 3.000 ;
        RECT  16.510 1.465 16.850 1.805 ;
        RECT  15.490 1.520 16.510 1.750 ;
        RECT  16.120 2.280 16.125 3.000 ;
        RECT  15.895 2.170 16.120 3.000 ;
        RECT  15.780 2.170 15.895 2.510 ;
        RECT  15.260 0.805 15.490 2.505 ;
        RECT  14.970 0.805 15.260 1.035 ;
        RECT  14.560 2.275 15.260 2.505 ;
        RECT  14.560 1.280 14.790 1.620 ;
        RECT  14.485 3.095 14.715 3.655 ;
        RECT  14.450 1.280 14.560 2.035 ;
        RECT  14.330 2.275 14.560 2.850 ;
        RECT  14.100 3.095 14.485 3.325 ;
        RECT  14.330 1.390 14.450 2.035 ;
        RECT  14.095 1.805 14.330 2.035 ;
        RECT  13.985 3.615 14.215 4.175 ;
        RECT  14.095 2.565 14.100 3.325 ;
        RECT  13.870 1.805 14.095 3.325 ;
        RECT  13.635 3.615 13.985 3.845 ;
        RECT  13.865 1.805 13.870 2.795 ;
        RECT  11.585 2.565 13.865 2.795 ;
        RECT  13.175 4.135 13.685 4.365 ;
        RECT  13.405 3.085 13.635 3.845 ;
        RECT  11.110 3.085 13.405 3.315 ;
        RECT  12.945 3.710 13.175 4.365 ;
        RECT  3.620 3.710 12.945 3.940 ;
        RECT  11.585 1.080 11.925 1.420 ;
        RECT  11.355 1.135 11.585 2.795 ;
        RECT  10.990 2.710 11.110 3.315 ;
        RECT  10.990 1.140 11.075 1.480 ;
        RECT  10.760 1.140 10.990 3.315 ;
        RECT  10.735 1.140 10.760 1.480 ;
        RECT  10.340 2.710 10.390 3.050 ;
        RECT  10.340 1.140 10.355 1.480 ;
        RECT  10.280 1.140 10.340 3.050 ;
        RECT  10.110 1.140 10.280 3.315 ;
        RECT  10.015 1.140 10.110 1.480 ;
        RECT  10.050 2.710 10.110 3.315 ;
        RECT  7.250 3.085 10.050 3.315 ;
        RECT  9.595 1.915 9.750 2.280 ;
        RECT  9.595 1.170 9.650 1.510 ;
        RECT  9.365 1.170 9.595 2.795 ;
        RECT  9.310 1.170 9.365 1.510 ;
        RECT  9.155 2.565 9.365 2.795 ;
        RECT  8.910 1.910 9.130 2.250 ;
        RECT  8.790 1.910 8.910 2.795 ;
        RECT  8.680 1.965 8.790 2.795 ;
        RECT  7.720 2.565 8.680 2.795 ;
        RECT  7.720 1.230 8.040 1.570 ;
        RECT  7.700 1.230 7.720 2.795 ;
        RECT  7.490 1.285 7.700 2.795 ;
        RECT  7.050 1.120 7.250 3.315 ;
        RECT  7.020 1.120 7.050 3.480 ;
        RECT  6.820 2.690 7.020 3.480 ;
        RECT  4.325 3.250 6.820 3.480 ;
        RECT  6.440 1.130 6.585 2.855 ;
        RECT  6.355 1.130 6.440 2.910 ;
        RECT  6.245 1.130 6.355 1.360 ;
        RECT  6.100 2.570 6.355 2.910 ;
        RECT  4.985 1.090 5.220 1.430 ;
        RECT  2.345 4.170 5.145 4.400 ;
        RECT  4.985 2.685 5.110 2.915 ;
        RECT  4.880 1.090 4.985 2.915 ;
        RECT  4.755 1.145 4.880 2.915 ;
        RECT  4.750 2.070 4.755 2.915 ;
        RECT  4.315 2.070 4.750 2.415 ;
        RECT  4.180 1.070 4.520 1.445 ;
        RECT  4.085 2.910 4.325 3.480 ;
        RECT  4.085 1.215 4.180 1.445 ;
        RECT  4.040 1.215 4.085 3.480 ;
        RECT  3.855 1.215 4.040 3.315 ;
        RECT  3.620 0.735 3.750 0.965 ;
        RECT  3.390 0.735 3.620 3.940 ;
        RECT  3.320 2.760 3.390 3.115 ;
        RECT  2.770 3.350 3.110 3.690 ;
        RECT  2.990 1.420 3.100 1.760 ;
        RECT  2.885 1.420 2.990 3.045 ;
        RECT  2.760 1.420 2.885 3.100 ;
        RECT  2.300 3.350 2.770 3.580 ;
        RECT  2.545 2.760 2.760 3.100 ;
        RECT  2.115 3.945 2.345 4.400 ;
        RECT  2.070 1.545 2.300 3.580 ;
        RECT  0.520 3.945 2.115 4.175 ;
        RECT  1.640 1.545 2.070 1.775 ;
        RECT  1.080 2.935 2.070 3.165 ;
        RECT  1.410 1.410 1.640 1.775 ;
        RECT  1.330 0.675 1.480 0.905 ;
        RECT  1.100 0.675 1.330 1.095 ;
        RECT  0.410 0.865 1.100 1.095 ;
        RECT  0.795 2.760 1.080 3.165 ;
        RECT  0.740 2.760 0.795 3.100 ;
        RECT  0.410 3.670 0.520 4.175 ;
        RECT  0.180 0.865 0.410 4.175 ;
    END
END SEDFFTRX1

MACRO SEDFFXL
    CLASS CORE ;
    FOREIGN SEDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 2.240 3.310 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 2.280 1.765 2.730 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.375 1.590 17.605 3.460 ;
        RECT  17.130 1.590 17.375 1.820 ;
        RECT  17.080 3.120 17.375 3.460 ;
        RECT  16.790 1.350 17.130 1.820 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.305 0.895 16.535 3.745 ;
        RECT  16.055 0.895 16.305 1.125 ;
        RECT  16.285 3.515 16.305 3.745 ;
        RECT  16.055 3.515 16.285 3.780 ;
        RECT  15.825 0.700 16.055 1.125 ;
        RECT  15.940 3.550 16.055 3.780 ;
        RECT  15.710 3.550 15.940 4.225 ;
        RECT  15.485 0.680 15.825 1.125 ;
        RECT  15.600 3.885 15.710 4.225 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.525 1.105 3.820 ;
        RECT  0.705 3.590 0.875 3.820 ;
        RECT  0.475 3.590 0.705 4.120 ;
        RECT  0.365 3.780 0.475 4.120 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 2.200 4.480 2.635 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.290 1.820 9.760 2.275 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.045 -0.400 17.820 0.400 ;
        RECT  16.705 -0.400 17.045 0.575 ;
        RECT  14.990 -0.400 16.705 0.400 ;
        RECT  14.760 -0.400 14.990 1.565 ;
        RECT  12.245 -0.400 14.760 0.400 ;
        RECT  11.905 -0.400 12.245 0.980 ;
        RECT  10.485 -0.400 11.905 0.400 ;
        RECT  10.145 -0.400 10.485 0.870 ;
        RECT  3.250 -0.400 10.145 0.400 ;
        RECT  3.020 -0.400 3.250 0.900 ;
        RECT  0.660 -0.400 3.020 0.400 ;
        RECT  0.320 -0.400 0.660 0.575 ;
        RECT  0.000 -0.400 0.320 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.200 4.640 17.820 5.440 ;
        RECT  16.805 4.465 17.200 5.440 ;
        RECT  15.175 4.610 16.805 5.440 ;
        RECT  14.835 3.400 15.175 5.440 ;
        RECT  12.495 4.640 14.835 5.440 ;
        RECT  11.555 4.465 12.495 5.440 ;
        RECT  10.460 4.640 11.555 5.440 ;
        RECT  8.960 4.465 10.460 5.440 ;
        RECT  2.950 4.640 8.960 5.440 ;
        RECT  2.610 3.980 2.950 5.440 ;
        RECT  1.410 4.640 2.610 5.440 ;
        RECT  1.070 4.080 1.410 5.440 ;
        RECT  0.000 4.640 1.070 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.945 1.515 16.075 3.185 ;
        RECT  15.865 1.515 15.945 3.240 ;
        RECT  15.845 1.460 15.865 3.240 ;
        RECT  15.525 1.460 15.845 1.800 ;
        RECT  15.605 2.885 15.845 3.240 ;
        RECT  14.760 2.885 15.605 3.115 ;
        RECT  14.470 2.100 15.460 2.440 ;
        RECT  14.420 2.830 14.760 3.170 ;
        RECT  14.240 0.685 14.470 2.440 ;
        RECT  14.375 2.940 14.420 3.170 ;
        RECT  14.145 2.940 14.375 4.175 ;
        RECT  13.280 0.685 14.240 0.915 ;
        RECT  13.910 2.210 14.240 2.440 ;
        RECT  6.770 3.945 14.145 4.175 ;
        RECT  13.450 1.255 14.010 1.485 ;
        RECT  13.755 2.210 13.910 3.425 ;
        RECT  13.680 2.210 13.755 3.590 ;
        RECT  13.525 3.195 13.680 3.590 ;
        RECT  13.290 1.255 13.450 2.765 ;
        RECT  13.220 1.255 13.290 3.655 ;
        RECT  13.060 2.535 13.220 3.655 ;
        RECT  9.800 3.425 13.060 3.655 ;
        RECT  12.600 1.415 12.830 3.135 ;
        RECT  11.610 1.415 12.600 1.645 ;
        RECT  11.580 2.905 12.600 3.135 ;
        RECT  12.030 2.290 12.370 2.630 ;
        RECT  11.120 2.345 12.030 2.575 ;
        RECT  11.270 0.675 11.610 1.680 ;
        RECT  10.715 0.675 11.270 0.905 ;
        RECT  10.855 2.345 11.120 3.100 ;
        RECT  10.710 1.280 10.855 3.100 ;
        RECT  10.625 1.280 10.710 3.030 ;
        RECT  8.855 2.800 10.625 3.030 ;
        RECT  10.165 1.315 10.395 2.155 ;
        RECT  9.915 1.315 10.165 1.545 ;
        RECT  9.685 0.675 9.915 1.545 ;
        RECT  9.460 3.260 9.800 3.655 ;
        RECT  8.255 0.675 9.685 0.905 ;
        RECT  8.395 3.425 9.460 3.655 ;
        RECT  9.200 1.250 9.430 1.590 ;
        RECT  8.395 1.360 9.200 1.590 ;
        RECT  8.625 2.145 8.855 3.030 ;
        RECT  8.165 1.360 8.395 3.655 ;
        RECT  8.025 0.675 8.255 1.110 ;
        RECT  6.965 1.885 8.165 2.115 ;
        RECT  8.010 3.425 8.165 3.655 ;
        RECT  7.625 0.880 8.025 1.110 ;
        RECT  7.825 2.840 7.935 3.180 ;
        RECT  7.595 2.380 7.825 3.180 ;
        RECT  7.515 0.880 7.625 1.220 ;
        RECT  6.660 2.380 7.595 2.610 ;
        RECT  7.285 0.880 7.515 1.645 ;
        RECT  6.660 1.415 7.285 1.645 ;
        RECT  6.795 2.840 7.135 3.180 ;
        RECT  6.575 0.955 6.825 1.185 ;
        RECT  6.195 2.950 6.795 3.180 ;
        RECT  6.540 3.500 6.770 4.175 ;
        RECT  6.430 1.415 6.660 2.610 ;
        RECT  6.345 0.685 6.575 1.185 ;
        RECT  6.430 3.500 6.540 3.840 ;
        RECT  3.895 0.685 6.345 0.915 ;
        RECT  5.965 2.950 6.195 4.410 ;
        RECT  4.620 4.180 5.965 4.410 ;
        RECT  5.390 3.505 5.730 3.950 ;
        RECT  5.360 1.735 5.690 2.160 ;
        RECT  2.790 1.250 5.465 1.480 ;
        RECT  2.380 3.505 5.390 3.735 ;
        RECT  5.130 1.735 5.360 3.275 ;
        RECT  2.325 1.735 5.130 1.965 ;
        RECT  4.925 3.045 5.130 3.275 ;
        RECT  4.390 4.015 4.620 4.410 ;
        RECT  3.970 4.015 4.390 4.245 ;
        RECT  3.565 2.920 3.905 3.260 ;
        RECT  2.410 2.975 3.565 3.205 ;
        RECT  2.560 0.630 2.790 1.480 ;
        RECT  1.730 0.630 2.560 0.860 ;
        RECT  2.070 2.310 2.410 3.205 ;
        RECT  2.150 3.505 2.380 4.110 ;
        RECT  2.095 1.090 2.325 1.965 ;
        RECT  1.810 3.770 2.150 4.110 ;
        RECT  0.520 1.090 2.095 1.320 ;
        RECT  1.920 2.975 2.070 3.205 ;
        RECT  1.690 2.975 1.920 3.310 ;
        RECT  1.635 1.580 1.865 1.960 ;
        RECT  0.995 2.975 1.690 3.205 ;
        RECT  0.995 1.730 1.635 1.960 ;
        RECT  0.765 1.730 0.995 3.205 ;
        RECT  0.465 1.090 0.520 1.780 ;
        RECT  0.465 2.970 0.520 3.310 ;
        RECT  0.290 1.090 0.465 3.310 ;
        RECT  0.235 1.440 0.290 3.310 ;
        RECT  0.180 1.440 0.235 1.780 ;
        RECT  0.180 2.970 0.235 3.310 ;
    END
END SEDFFXL

MACRO SEDFFX4
    CLASS CORE ;
    FOREIGN SEDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 2.220 3.945 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 2.280 1.985 2.635 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.640 1.395 22.215 1.735 ;
        RECT  21.620 2.900 22.050 3.240 ;
        RECT  21.620 1.260 21.640 2.660 ;
        RECT  21.280 1.260 21.620 3.240 ;
        RECT  21.260 1.260 21.280 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.960 1.260 20.980 2.660 ;
        RECT  20.620 1.260 20.960 3.240 ;
        RECT  20.600 1.260 20.620 2.660 ;
        RECT  20.430 2.900 20.620 3.240 ;
        RECT  20.595 1.390 20.600 1.730 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 3.525 1.105 3.755 ;
        RECT  0.775 3.525 1.005 4.010 ;
        RECT  0.740 3.780 0.775 4.010 ;
        RECT  0.400 3.780 0.740 4.120 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.950 2.405 5.065 2.635 ;
        RECT  4.555 2.405 4.950 2.915 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.740 1.820 10.420 2.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.920 -0.400 23.100 0.400 ;
        RECT  22.580 -0.400 22.920 1.100 ;
        RECT  21.575 -0.400 22.580 0.400 ;
        RECT  21.235 -0.400 21.575 0.990 ;
        RECT  20.290 -0.400 21.235 0.400 ;
        RECT  19.950 -0.400 20.290 0.955 ;
        RECT  18.870 -0.400 19.950 0.400 ;
        RECT  18.530 -0.400 18.870 1.680 ;
        RECT  16.115 -0.400 18.530 0.400 ;
        RECT  15.775 -0.400 16.115 0.575 ;
        RECT  13.515 -0.400 15.775 0.400 ;
        RECT  13.175 -0.400 13.515 1.010 ;
        RECT  11.140 -0.400 13.175 0.400 ;
        RECT  10.800 -0.400 11.140 1.000 ;
        RECT  3.415 -0.400 10.800 0.400 ;
        RECT  3.075 -0.400 3.415 0.970 ;
        RECT  0.640 -0.400 3.075 0.400 ;
        RECT  0.300 -0.400 0.640 0.575 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.730 4.640 23.100 5.440 ;
        RECT  22.390 3.990 22.730 5.440 ;
        RECT  21.410 4.640 22.390 5.440 ;
        RECT  21.070 4.090 21.410 5.440 ;
        RECT  20.130 4.640 21.070 5.440 ;
        RECT  19.790 4.090 20.130 5.440 ;
        RECT  18.650 4.640 19.790 5.440 ;
        RECT  18.220 4.465 18.650 5.440 ;
        RECT  15.820 4.640 18.220 5.440 ;
        RECT  15.480 4.465 15.820 5.440 ;
        RECT  12.965 4.640 15.480 5.440 ;
        RECT  12.625 4.465 12.965 5.440 ;
        RECT  10.705 4.640 12.625 5.440 ;
        RECT  10.365 4.465 10.705 5.440 ;
        RECT  9.400 4.640 10.365 5.440 ;
        RECT  9.060 4.465 9.400 5.440 ;
        RECT  3.270 4.640 9.060 5.440 ;
        RECT  2.930 3.890 3.270 5.440 ;
        RECT  1.750 4.640 2.930 5.440 ;
        RECT  1.410 3.800 1.750 5.440 ;
        RECT  0.000 4.640 1.410 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.510 2.200 22.685 2.540 ;
        RECT  22.280 2.200 22.510 3.700 ;
        RECT  21.875 2.200 22.280 2.540 ;
        RECT  20.015 3.470 22.280 3.700 ;
        RECT  19.785 1.435 20.015 3.700 ;
        RECT  19.590 1.435 19.785 1.665 ;
        RECT  19.410 3.390 19.785 3.700 ;
        RECT  19.250 0.855 19.590 1.665 ;
        RECT  18.835 3.390 19.410 3.730 ;
        RECT  18.375 1.980 19.345 2.320 ;
        RECT  18.605 2.690 18.835 4.175 ;
        RECT  14.995 3.945 18.605 4.175 ;
        RECT  18.290 1.980 18.375 3.655 ;
        RECT  18.145 1.055 18.290 3.655 ;
        RECT  18.060 1.055 18.145 2.210 ;
        RECT  14.445 3.425 18.145 3.655 ;
        RECT  17.435 1.055 18.060 1.285 ;
        RECT  17.510 1.645 17.740 2.955 ;
        RECT  16.425 2.725 17.510 2.955 ;
        RECT  17.095 0.945 17.435 1.285 ;
        RECT  14.795 0.945 17.095 1.175 ;
        RECT  16.810 1.615 17.040 1.980 ;
        RECT  13.525 1.615 16.810 1.845 ;
        RECT  16.085 2.115 16.425 2.955 ;
        RECT  13.985 2.725 16.085 2.955 ;
        RECT  14.765 3.945 14.995 4.410 ;
        RECT  14.455 0.835 14.795 1.175 ;
        RECT  13.580 4.180 14.765 4.410 ;
        RECT  14.215 3.425 14.445 3.950 ;
        RECT  13.755 2.725 13.985 3.655 ;
        RECT  8.365 3.425 13.755 3.655 ;
        RECT  13.350 4.005 13.580 4.410 ;
        RECT  13.295 1.335 13.525 3.075 ;
        RECT  8.735 4.005 13.350 4.235 ;
        RECT  12.755 1.335 13.295 1.565 ;
        RECT  11.860 2.845 13.295 3.075 ;
        RECT  12.830 2.120 13.060 2.550 ;
        RECT  11.630 2.120 12.830 2.350 ;
        RECT  12.455 1.200 12.755 1.565 ;
        RECT  12.225 0.685 12.455 1.565 ;
        RECT  12.055 0.685 12.225 0.915 ;
        RECT  11.630 1.210 11.810 1.710 ;
        RECT  11.580 1.210 11.630 3.055 ;
        RECT  11.400 1.480 11.580 3.055 ;
        RECT  8.945 2.825 11.400 3.055 ;
        RECT  10.940 1.315 11.170 2.330 ;
        RECT  10.570 1.315 10.940 1.545 ;
        RECT  10.340 0.630 10.570 1.545 ;
        RECT  8.185 0.630 10.340 0.860 ;
        RECT  9.770 1.220 10.110 1.560 ;
        RECT  9.135 1.330 9.770 1.560 ;
        RECT  8.905 1.330 9.135 1.835 ;
        RECT  8.715 2.270 8.945 3.055 ;
        RECT  8.365 1.605 8.905 1.835 ;
        RECT  8.505 4.005 8.735 4.365 ;
        RECT  6.665 4.135 8.505 4.365 ;
        RECT  8.135 1.605 8.365 3.720 ;
        RECT  8.075 0.630 8.185 1.240 ;
        RECT  7.410 1.605 8.135 1.835 ;
        RECT  7.990 3.490 8.135 3.720 ;
        RECT  7.955 0.630 8.075 1.375 ;
        RECT  7.845 0.900 7.955 1.375 ;
        RECT  7.700 2.595 7.905 3.245 ;
        RECT  7.145 1.145 7.845 1.375 ;
        RECT  7.675 2.255 7.700 3.245 ;
        RECT  7.470 2.255 7.675 2.825 ;
        RECT  7.145 2.255 7.470 2.485 ;
        RECT  5.990 0.685 7.420 0.915 ;
        RECT  6.900 3.100 7.240 3.440 ;
        RECT  6.915 1.145 7.145 2.485 ;
        RECT  6.425 3.210 6.900 3.440 ;
        RECT  6.195 3.210 6.425 4.225 ;
        RECT  5.600 1.775 6.340 2.005 ;
        RECT  4.640 3.995 6.195 4.225 ;
        RECT  2.840 1.205 6.100 1.435 ;
        RECT  5.760 0.685 5.990 0.970 ;
        RECT  5.245 3.505 5.960 3.735 ;
        RECT  4.435 0.740 5.760 0.970 ;
        RECT  5.370 1.725 5.600 3.165 ;
        RECT  2.380 1.725 5.370 1.955 ;
        RECT  5.250 2.935 5.370 3.165 ;
        RECT  5.015 3.425 5.245 3.735 ;
        RECT  2.510 3.425 5.015 3.655 ;
        RECT  4.300 3.885 4.640 4.225 ;
        RECT  2.865 2.890 4.225 3.120 ;
        RECT  2.865 2.185 2.920 2.525 ;
        RECT  2.635 2.185 2.865 3.195 ;
        RECT  2.610 0.695 2.840 1.435 ;
        RECT  2.580 2.185 2.635 2.525 ;
        RECT  1.970 2.965 2.635 3.195 ;
        RECT  2.080 0.695 2.610 0.925 ;
        RECT  2.280 3.425 2.510 4.110 ;
        RECT  2.150 1.155 2.380 1.955 ;
        RECT  2.170 3.770 2.280 4.110 ;
        RECT  0.520 1.155 2.150 1.385 ;
        RECT  1.630 2.965 1.970 3.360 ;
        RECT  1.065 1.615 1.920 1.845 ;
        RECT  1.065 2.965 1.630 3.195 ;
        RECT  0.835 1.615 1.065 3.195 ;
        RECT  0.465 1.155 0.520 1.780 ;
        RECT  0.290 1.155 0.465 3.360 ;
        RECT  0.235 1.440 0.290 3.360 ;
        RECT  0.180 1.440 0.235 1.780 ;
    END
END SEDFFX4

MACRO SEDFFX2
    CLASS CORE ;
    FOREIGN SEDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 2.240 3.330 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.420 2.185 1.895 2.695 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.390 1.285 19.620 4.030 ;
        RECT  19.355 1.285 19.390 1.705 ;
        RECT  19.280 3.090 19.390 4.030 ;
        RECT  19.240 1.365 19.355 1.705 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.265 1.365 18.295 1.845 ;
        RECT  18.240 1.285 18.265 1.845 ;
        RECT  18.120 1.285 18.240 2.965 ;
        RECT  18.010 1.285 18.120 3.200 ;
        RECT  17.960 1.365 18.010 1.845 ;
        RECT  17.890 2.540 18.010 3.200 ;
        RECT  17.955 1.365 17.960 1.705 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 3.525 1.105 3.755 ;
        RECT  0.750 3.525 0.925 4.010 ;
        RECT  0.695 3.525 0.750 4.120 ;
        RECT  0.410 3.780 0.695 4.120 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.915 2.255 4.480 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 1.820 9.795 2.370 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.940 -0.400 19.800 0.400 ;
        RECT  18.600 -0.400 18.940 0.990 ;
        RECT  16.935 -0.400 18.600 0.400 ;
        RECT  16.595 -0.400 16.935 1.400 ;
        RECT  14.935 -0.400 16.595 0.400 ;
        RECT  16.590 1.060 16.595 1.345 ;
        RECT  14.595 -0.400 14.935 1.060 ;
        RECT  12.290 -0.400 14.595 0.400 ;
        RECT  11.950 -0.400 12.290 0.860 ;
        RECT  10.510 -0.400 11.950 0.400 ;
        RECT  10.170 -0.400 10.510 0.900 ;
        RECT  3.410 -0.400 10.170 0.400 ;
        RECT  3.070 -0.400 3.410 0.815 ;
        RECT  0.640 -0.400 3.070 0.400 ;
        RECT  0.300 -0.400 0.640 0.575 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.900 4.640 19.800 5.440 ;
        RECT  18.560 4.075 18.900 5.440 ;
        RECT  16.715 4.630 18.560 5.440 ;
        RECT  15.215 4.465 16.715 5.440 ;
        RECT  12.455 4.640 15.215 5.440 ;
        RECT  11.435 4.465 12.455 5.440 ;
        RECT  10.115 4.640 11.435 5.440 ;
        RECT  8.835 4.465 10.115 5.440 ;
        RECT  2.955 4.640 8.835 5.440 ;
        RECT  2.615 3.895 2.955 5.440 ;
        RECT  1.495 4.640 2.615 5.440 ;
        RECT  1.155 4.010 1.495 5.440 ;
        RECT  0.000 4.640 1.155 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.965 2.160 19.160 2.695 ;
        RECT  18.930 2.160 18.965 3.845 ;
        RECT  18.735 2.465 18.930 3.845 ;
        RECT  17.475 3.615 18.735 3.845 ;
        RECT  17.475 1.170 17.540 2.885 ;
        RECT  17.310 1.170 17.475 3.965 ;
        RECT  17.245 2.655 17.310 3.965 ;
        RECT  17.135 3.080 17.245 3.965 ;
        RECT  16.715 3.735 17.135 3.965 ;
        RECT  16.740 1.850 16.970 2.215 ;
        RECT  16.255 1.855 16.740 2.215 ;
        RECT  16.485 3.735 16.715 4.030 ;
        RECT  16.250 3.800 16.485 4.030 ;
        RECT  16.025 1.555 16.255 3.010 ;
        RECT  15.910 3.800 16.250 4.235 ;
        RECT  15.515 1.555 16.025 1.785 ;
        RECT  15.855 2.780 16.025 3.010 ;
        RECT  8.605 4.005 15.910 4.235 ;
        RECT  15.515 2.780 15.855 3.120 ;
        RECT  15.455 2.100 15.795 2.440 ;
        RECT  15.175 1.420 15.515 1.785 ;
        RECT  14.735 2.890 15.515 3.120 ;
        RECT  14.105 2.210 15.455 2.440 ;
        RECT  14.105 1.555 15.175 1.785 ;
        RECT  14.505 2.890 14.735 3.520 ;
        RECT  13.855 3.290 14.505 3.520 ;
        RECT  13.875 1.240 14.105 1.785 ;
        RECT  13.875 2.210 14.105 2.765 ;
        RECT  13.610 1.240 13.875 1.470 ;
        RECT  13.485 2.535 13.875 2.765 ;
        RECT  13.515 3.290 13.855 3.630 ;
        RECT  13.270 1.130 13.610 1.470 ;
        RECT  12.370 1.855 13.600 2.085 ;
        RECT  13.145 2.535 13.485 2.890 ;
        RECT  13.050 2.660 13.145 2.890 ;
        RECT  12.820 2.660 13.050 3.670 ;
        RECT  9.610 3.440 12.820 3.670 ;
        RECT  12.140 1.415 12.370 3.210 ;
        RECT  11.690 1.415 12.140 1.645 ;
        RECT  11.535 2.980 12.140 3.210 ;
        RECT  10.930 2.455 11.905 2.685 ;
        RECT  11.580 1.280 11.690 1.645 ;
        RECT  11.405 0.675 11.580 1.645 ;
        RECT  11.350 0.675 11.405 1.620 ;
        RECT  10.835 0.675 11.350 0.905 ;
        RECT  10.700 1.400 10.930 3.075 ;
        RECT  10.485 2.815 10.700 3.075 ;
        RECT  8.595 2.815 10.485 3.045 ;
        RECT  10.185 1.315 10.415 2.310 ;
        RECT  9.940 1.315 10.185 1.545 ;
        RECT  9.710 0.675 9.940 1.545 ;
        RECT  8.475 0.675 9.710 0.905 ;
        RECT  9.215 3.285 9.610 3.670 ;
        RECT  9.200 1.190 9.430 1.590 ;
        RECT  8.135 3.285 9.215 3.515 ;
        RECT  9.150 1.360 9.200 1.590 ;
        RECT  8.920 1.360 9.150 1.865 ;
        RECT  8.135 1.635 8.920 1.865 ;
        RECT  8.375 4.005 8.605 4.410 ;
        RECT  8.365 2.180 8.595 3.045 ;
        RECT  8.245 0.675 8.475 1.105 ;
        RECT  6.710 4.180 8.375 4.410 ;
        RECT  7.625 0.875 8.245 1.105 ;
        RECT  7.905 1.635 8.135 3.830 ;
        RECT  6.865 1.645 7.905 1.875 ;
        RECT  7.755 3.600 7.905 3.830 ;
        RECT  7.440 2.255 7.670 3.280 ;
        RECT  7.515 0.875 7.625 1.260 ;
        RECT  7.285 0.875 7.515 1.410 ;
        RECT  6.400 2.255 7.440 2.485 ;
        RECT  6.400 1.180 7.285 1.410 ;
        RECT  6.665 2.940 7.005 3.280 ;
        RECT  3.960 0.655 6.825 0.885 ;
        RECT  6.480 3.950 6.710 4.410 ;
        RECT  6.145 3.050 6.665 3.280 ;
        RECT  6.170 1.180 6.400 2.485 ;
        RECT  5.915 3.050 6.145 4.395 ;
        RECT  4.450 4.165 5.915 4.395 ;
        RECT  5.315 1.695 5.870 1.925 ;
        RECT  5.310 3.705 5.685 3.935 ;
        RECT  5.350 1.165 5.460 1.395 ;
        RECT  5.120 1.115 5.350 1.395 ;
        RECT  5.085 1.695 5.315 3.200 ;
        RECT  5.080 3.435 5.310 3.935 ;
        RECT  2.840 1.115 5.120 1.345 ;
        RECT  4.760 1.695 5.085 1.925 ;
        RECT  4.930 2.970 5.085 3.200 ;
        RECT  2.385 3.435 5.080 3.665 ;
        RECT  4.530 1.575 4.760 1.925 ;
        RECT  2.380 1.575 4.530 1.805 ;
        RECT  4.220 3.900 4.450 4.395 ;
        RECT  3.975 3.900 4.220 4.130 ;
        RECT  2.380 2.975 3.905 3.205 ;
        RECT  2.610 0.690 2.840 1.345 ;
        RECT  1.880 0.690 2.610 0.920 ;
        RECT  2.380 2.035 2.530 2.265 ;
        RECT  2.195 3.435 2.385 4.000 ;
        RECT  2.150 1.150 2.380 1.805 ;
        RECT  2.150 2.035 2.380 3.205 ;
        RECT  2.155 3.435 2.195 4.110 ;
        RECT  1.855 3.770 2.155 4.110 ;
        RECT  0.520 1.150 2.150 1.380 ;
        RECT  1.880 2.930 2.150 3.205 ;
        RECT  1.155 1.610 1.920 1.840 ;
        RECT  1.540 2.930 1.880 3.270 ;
        RECT  1.155 2.930 1.540 3.160 ;
        RECT  0.925 1.610 1.155 3.160 ;
        RECT  0.465 1.150 0.520 1.780 ;
        RECT  0.290 1.150 0.465 3.360 ;
        RECT  0.235 1.440 0.290 3.360 ;
        RECT  0.180 1.440 0.235 1.780 ;
    END
END SEDFFX2

MACRO SEDFFX1
    CLASS CORE ;
    FOREIGN SEDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 2.240 3.310 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 2.280 1.765 2.730 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.375 1.590 17.605 3.460 ;
        RECT  17.130 1.590 17.375 1.820 ;
        RECT  17.080 3.120 17.375 3.460 ;
        RECT  16.790 1.345 17.130 1.820 ;
        RECT  16.785 1.400 16.790 1.820 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.305 0.895 16.535 3.745 ;
        RECT  16.055 0.895 16.305 1.125 ;
        RECT  16.285 3.515 16.305 3.745 ;
        RECT  16.055 3.515 16.285 3.780 ;
        RECT  15.485 0.735 16.055 1.125 ;
        RECT  15.940 3.550 16.055 3.780 ;
        RECT  15.710 3.550 15.940 4.225 ;
        RECT  15.600 3.885 15.710 4.225 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.525 1.105 3.820 ;
        RECT  0.705 3.590 0.875 3.820 ;
        RECT  0.475 3.590 0.705 4.120 ;
        RECT  0.365 3.780 0.475 4.120 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 2.200 4.480 2.635 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.290 1.820 9.760 2.275 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.045 -0.400 17.820 0.400 ;
        RECT  16.705 -0.400 17.045 0.575 ;
        RECT  14.990 -0.400 16.705 0.400 ;
        RECT  14.760 -0.400 14.990 1.495 ;
        RECT  12.245 -0.400 14.760 0.400 ;
        RECT  11.905 -0.400 12.245 0.980 ;
        RECT  10.485 -0.400 11.905 0.400 ;
        RECT  10.145 -0.400 10.485 0.870 ;
        RECT  3.250 -0.400 10.145 0.400 ;
        RECT  3.020 -0.400 3.250 0.900 ;
        RECT  0.660 -0.400 3.020 0.400 ;
        RECT  0.320 -0.400 0.660 0.575 ;
        RECT  0.000 -0.400 0.320 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.200 4.640 17.820 5.440 ;
        RECT  16.805 4.465 17.200 5.440 ;
        RECT  15.175 4.610 16.805 5.440 ;
        RECT  14.835 3.490 15.175 5.440 ;
        RECT  12.490 4.640 14.835 5.440 ;
        RECT  11.550 4.465 12.490 5.440 ;
        RECT  10.460 4.640 11.550 5.440 ;
        RECT  8.960 4.465 10.460 5.440 ;
        RECT  2.950 4.640 8.960 5.440 ;
        RECT  2.610 3.980 2.950 5.440 ;
        RECT  1.410 4.640 2.610 5.440 ;
        RECT  1.070 4.080 1.410 5.440 ;
        RECT  0.000 4.640 1.070 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.865 1.515 16.075 3.160 ;
        RECT  15.845 1.460 15.865 3.160 ;
        RECT  15.525 1.460 15.845 1.800 ;
        RECT  15.605 2.820 15.845 3.160 ;
        RECT  14.760 2.895 15.605 3.125 ;
        RECT  14.470 2.100 15.460 2.440 ;
        RECT  14.420 2.840 14.760 3.180 ;
        RECT  14.240 0.685 14.470 2.440 ;
        RECT  14.375 2.950 14.420 3.180 ;
        RECT  14.145 2.950 14.375 4.175 ;
        RECT  13.280 0.685 14.240 0.915 ;
        RECT  13.910 2.210 14.240 2.440 ;
        RECT  6.770 3.945 14.145 4.175 ;
        RECT  13.450 1.255 14.010 1.485 ;
        RECT  13.680 2.210 13.910 3.425 ;
        RECT  13.525 3.060 13.680 3.425 ;
        RECT  13.290 1.255 13.450 2.765 ;
        RECT  13.220 1.255 13.290 3.655 ;
        RECT  13.060 2.535 13.220 3.655 ;
        RECT  11.255 3.425 13.060 3.655 ;
        RECT  12.600 1.415 12.830 3.135 ;
        RECT  11.610 1.415 12.600 1.645 ;
        RECT  11.580 2.905 12.600 3.135 ;
        RECT  12.030 2.290 12.370 2.630 ;
        RECT  11.120 2.345 12.030 2.575 ;
        RECT  11.270 0.675 11.610 1.680 ;
        RECT  10.715 0.675 11.270 0.905 ;
        RECT  9.800 3.385 11.255 3.655 ;
        RECT  10.855 2.345 11.120 3.100 ;
        RECT  10.835 1.280 10.855 3.100 ;
        RECT  10.625 1.280 10.835 2.575 ;
        RECT  8.855 2.870 10.835 3.100 ;
        RECT  10.165 1.315 10.395 2.155 ;
        RECT  9.915 1.315 10.165 1.545 ;
        RECT  9.685 0.675 9.915 1.545 ;
        RECT  9.460 3.330 9.800 3.670 ;
        RECT  8.255 0.675 9.685 0.905 ;
        RECT  8.395 3.425 9.460 3.655 ;
        RECT  9.200 1.250 9.430 1.590 ;
        RECT  8.395 1.360 9.200 1.590 ;
        RECT  8.625 2.145 8.855 3.100 ;
        RECT  8.165 1.360 8.395 3.655 ;
        RECT  8.025 0.675 8.255 1.110 ;
        RECT  6.965 1.885 8.165 2.115 ;
        RECT  8.010 3.425 8.165 3.655 ;
        RECT  7.625 0.880 8.025 1.110 ;
        RECT  7.825 2.840 7.935 3.180 ;
        RECT  7.595 2.380 7.825 3.180 ;
        RECT  7.515 0.880 7.625 1.220 ;
        RECT  6.660 2.380 7.595 2.610 ;
        RECT  7.285 0.880 7.515 1.645 ;
        RECT  6.660 1.415 7.285 1.645 ;
        RECT  6.795 2.840 7.135 3.180 ;
        RECT  6.575 0.955 6.825 1.185 ;
        RECT  6.195 2.950 6.795 3.180 ;
        RECT  6.540 3.500 6.770 4.175 ;
        RECT  6.430 1.415 6.660 2.610 ;
        RECT  6.345 0.685 6.575 1.185 ;
        RECT  6.430 3.500 6.540 3.840 ;
        RECT  3.895 0.685 6.345 0.915 ;
        RECT  5.965 2.950 6.195 4.410 ;
        RECT  4.620 4.180 5.965 4.410 ;
        RECT  5.390 3.505 5.730 3.950 ;
        RECT  5.360 1.735 5.690 2.160 ;
        RECT  2.790 1.250 5.465 1.480 ;
        RECT  2.380 3.505 5.390 3.735 ;
        RECT  5.130 1.735 5.360 3.275 ;
        RECT  2.325 1.735 5.130 1.965 ;
        RECT  4.925 3.045 5.130 3.275 ;
        RECT  4.390 4.015 4.620 4.410 ;
        RECT  3.970 4.015 4.390 4.245 ;
        RECT  3.565 2.920 3.905 3.260 ;
        RECT  2.410 2.975 3.565 3.205 ;
        RECT  2.560 0.630 2.790 1.480 ;
        RECT  1.730 0.630 2.560 0.860 ;
        RECT  2.070 2.310 2.410 3.205 ;
        RECT  2.150 3.505 2.380 4.135 ;
        RECT  2.095 1.090 2.325 1.965 ;
        RECT  1.810 3.870 2.150 4.210 ;
        RECT  0.520 1.090 2.095 1.320 ;
        RECT  1.920 2.975 2.070 3.205 ;
        RECT  1.690 2.975 1.920 3.360 ;
        RECT  1.635 1.580 1.865 1.960 ;
        RECT  0.995 2.975 1.690 3.205 ;
        RECT  0.995 1.730 1.635 1.960 ;
        RECT  0.765 1.730 0.995 3.205 ;
        RECT  0.465 1.090 0.520 1.780 ;
        RECT  0.465 3.020 0.520 3.360 ;
        RECT  0.290 1.090 0.465 3.360 ;
        RECT  0.235 1.440 0.290 3.360 ;
        RECT  0.180 1.440 0.235 1.780 ;
        RECT  0.180 3.020 0.235 3.360 ;
    END
END SEDFFX1

MACRO SEDFFHQXL
    CLASS CORE ;
    FOREIGN SEDFFHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 0.685 1.945 1.085 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.060 1.105 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.015 1.360 20.245 3.240 ;
        RECT  19.830 1.360 20.015 1.700 ;
        RECT  19.895 2.900 20.015 3.240 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 2.275 7.120 2.630 ;
        RECT  6.815 2.275 7.045 2.635 ;
        RECT  6.430 2.275 6.815 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 0.725 5.065 1.040 ;
        RECT  4.415 0.810 4.835 1.040 ;
        RECT  4.415 2.005 4.435 2.370 ;
        RECT  4.205 0.810 4.415 2.370 ;
        RECT  4.185 0.810 4.205 2.235 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.310 1.770 9.995 2.150 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.610 -0.400 20.460 0.400 ;
        RECT  19.270 -0.400 19.610 0.575 ;
        RECT  18.475 -0.400 19.270 0.400 ;
        RECT  18.135 -0.400 18.475 0.575 ;
        RECT  15.270 -0.400 18.135 0.400 ;
        RECT  14.930 -0.400 15.270 1.595 ;
        RECT  12.965 -0.400 14.930 0.400 ;
        RECT  12.625 -0.400 12.965 1.270 ;
        RECT  10.410 -0.400 12.625 0.400 ;
        RECT  10.070 -0.400 10.410 0.575 ;
        RECT  7.045 -0.400 10.070 0.400 ;
        RECT  6.705 -0.400 7.045 0.575 ;
        RECT  4.345 -0.400 6.705 0.400 ;
        RECT  4.005 -0.400 4.345 0.575 ;
        RECT  1.120 -0.400 4.005 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.185 4.640 20.460 5.440 ;
        RECT  19.745 4.465 20.185 5.440 ;
        RECT  18.210 4.640 19.745 5.440 ;
        RECT  17.870 4.465 18.210 5.440 ;
        RECT  12.315 4.640 17.870 5.440 ;
        RECT  11.975 4.465 12.315 5.440 ;
        RECT  10.210 4.640 11.975 5.440 ;
        RECT  9.980 3.720 10.210 5.440 ;
        RECT  6.910 4.640 9.980 5.440 ;
        RECT  6.570 4.465 6.910 5.440 ;
        RECT  4.225 4.640 6.570 5.440 ;
        RECT  3.885 4.465 4.225 5.440 ;
        RECT  1.180 4.640 3.885 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.415 2.100 19.755 2.440 ;
        RECT  18.920 2.155 19.415 2.385 ;
        RECT  18.920 3.420 18.975 3.760 ;
        RECT  18.910 1.345 18.920 3.820 ;
        RECT  18.690 1.290 18.910 3.820 ;
        RECT  18.570 1.290 18.690 1.630 ;
        RECT  18.635 3.420 18.690 3.820 ;
        RECT  17.835 3.590 18.635 3.820 ;
        RECT  18.120 2.200 18.460 2.540 ;
        RECT  17.770 2.200 18.120 2.430 ;
        RECT  17.835 2.870 17.890 3.210 ;
        RECT  17.605 2.870 17.835 3.820 ;
        RECT  17.540 0.695 17.770 2.430 ;
        RECT  17.550 2.870 17.605 3.210 ;
        RECT  16.880 3.590 17.605 3.820 ;
        RECT  16.775 0.695 17.540 0.925 ;
        RECT  17.095 2.200 17.540 2.430 ;
        RECT  17.075 1.245 17.305 1.625 ;
        RECT  16.880 2.200 17.095 3.240 ;
        RECT  16.480 1.395 17.075 1.625 ;
        RECT  16.865 2.200 16.880 3.360 ;
        RECT  16.650 3.590 16.880 4.410 ;
        RECT  16.650 3.010 16.865 3.360 ;
        RECT  16.545 0.695 16.775 1.165 ;
        RECT  12.780 4.180 16.650 4.410 ;
        RECT  16.420 1.395 16.480 2.735 ;
        RECT  16.250 1.395 16.420 3.950 ;
        RECT  16.210 2.350 16.250 3.950 ;
        RECT  16.190 2.505 16.210 3.950 ;
        RECT  13.245 3.720 16.190 3.950 ;
        RECT  15.960 1.255 16.015 1.960 ;
        RECT  15.785 1.255 15.960 3.220 ;
        RECT  15.730 1.730 15.785 3.220 ;
        RECT  15.250 2.135 15.480 3.490 ;
        RECT  13.710 3.260 15.250 3.490 ;
        RECT  14.245 2.800 14.565 3.030 ;
        RECT  14.245 1.330 14.470 1.560 ;
        RECT  14.015 0.630 14.245 3.030 ;
        RECT  13.480 0.980 13.710 3.490 ;
        RECT  12.295 2.325 13.480 2.555 ;
        RECT  13.015 3.540 13.245 3.950 ;
        RECT  11.755 1.590 13.230 1.940 ;
        RECT  11.130 3.540 13.015 3.770 ;
        RECT  12.550 4.005 12.780 4.410 ;
        RECT  10.670 4.005 12.550 4.235 ;
        RECT  11.590 1.025 11.755 2.730 ;
        RECT  11.525 1.025 11.590 3.290 ;
        RECT  11.265 1.025 11.525 1.255 ;
        RECT  11.360 2.500 11.525 3.290 ;
        RECT  10.455 1.655 11.235 1.885 ;
        RECT  10.900 2.795 11.130 3.770 ;
        RECT  10.455 2.795 10.900 3.025 ;
        RECT  10.440 3.260 10.670 4.235 ;
        RECT  10.225 1.080 10.455 3.025 ;
        RECT  8.930 3.260 10.440 3.490 ;
        RECT  9.735 1.080 10.225 1.310 ;
        RECT  9.165 2.795 10.225 3.025 ;
        RECT  9.505 0.675 9.735 1.310 ;
        RECT  9.265 0.675 9.505 0.905 ;
        RECT  7.500 4.125 9.325 4.355 ;
        RECT  8.930 1.460 8.945 2.020 ;
        RECT  8.905 1.460 8.930 3.790 ;
        RECT  8.715 1.460 8.905 3.845 ;
        RECT  8.700 1.790 8.715 3.845 ;
        RECT  8.675 3.260 8.700 3.845 ;
        RECT  8.220 1.640 8.390 3.810 ;
        RECT  8.160 1.390 8.220 3.810 ;
        RECT  7.990 1.390 8.160 1.870 ;
        RECT  7.895 3.500 8.160 3.810 ;
        RECT  7.760 2.275 7.930 2.650 ;
        RECT  7.790 0.630 7.925 0.860 ;
        RECT  5.500 3.500 7.895 3.730 ;
        RECT  7.760 0.630 7.790 1.035 ;
        RECT  7.615 0.630 7.760 2.650 ;
        RECT  7.530 0.630 7.615 3.165 ;
        RECT  6.250 0.805 7.530 1.035 ;
        RECT  7.385 2.420 7.530 3.165 ;
        RECT  7.270 4.005 7.500 4.355 ;
        RECT  7.070 1.540 7.300 1.915 ;
        RECT  2.545 4.005 7.270 4.235 ;
        RECT  6.395 1.540 7.070 1.770 ;
        RECT  6.130 1.265 6.395 1.770 ;
        RECT  6.130 2.860 6.295 3.090 ;
        RECT  6.020 0.655 6.250 1.035 ;
        RECT  6.025 1.265 6.130 3.090 ;
        RECT  5.900 1.540 6.025 3.090 ;
        RECT  5.445 0.655 6.020 0.885 ;
        RECT  5.690 2.145 5.900 2.490 ;
        RECT  5.455 1.205 5.615 1.725 ;
        RECT  5.455 2.765 5.500 3.730 ;
        RECT  5.385 1.205 5.455 3.730 ;
        RECT  5.270 1.495 5.385 3.730 ;
        RECT  5.225 1.495 5.270 2.995 ;
        RECT  3.950 3.500 5.270 3.730 ;
        RECT  4.890 1.545 4.950 3.150 ;
        RECT  4.720 1.275 4.890 3.150 ;
        RECT  4.660 1.275 4.720 1.775 ;
        RECT  4.495 2.920 4.720 3.150 ;
        RECT  3.720 0.850 3.950 3.730 ;
        RECT  3.500 0.850 3.720 1.080 ;
        RECT  3.030 3.500 3.720 3.730 ;
        RECT  3.270 0.685 3.500 1.080 ;
        RECT  3.255 1.395 3.485 2.965 ;
        RECT  3.150 0.685 3.270 0.915 ;
        RECT  3.135 2.150 3.255 2.965 ;
        RECT  2.605 2.570 3.135 2.965 ;
        RECT  2.435 1.320 2.665 2.175 ;
        RECT  2.375 3.445 2.545 4.235 ;
        RECT  2.375 1.945 2.435 2.175 ;
        RECT  2.315 1.945 2.375 4.235 ;
        RECT  2.145 1.945 2.315 3.730 ;
        RECT  1.680 4.140 2.085 4.370 ;
        RECT  1.810 1.455 1.920 1.685 ;
        RECT  1.810 3.135 1.840 3.475 ;
        RECT  1.580 1.455 1.810 3.475 ;
        RECT  1.450 3.770 1.680 4.370 ;
        RECT  1.500 3.135 1.580 3.475 ;
        RECT  0.520 3.770 1.450 4.000 ;
        RECT  0.410 1.440 0.520 1.780 ;
        RECT  0.410 3.135 0.520 4.000 ;
        RECT  0.290 1.440 0.410 4.000 ;
        RECT  0.180 1.440 0.290 3.475 ;
    END
END SEDFFHQXL

MACRO SEDFFHQX4
    CLASS CORE ;
    FOREIGN SEDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFHQXL ;
    SIZE 25.080 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 0.700 1.945 1.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.060 1.105 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.075 1.820 24.280 3.220 ;
        RECT  23.900 1.450 24.075 3.220 ;
        RECT  23.735 1.450 23.900 3.080 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.740 2.305 7.120 2.910 ;
        RECT  6.475 2.330 6.740 2.560 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.485 2.370 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 2.075 9.900 2.415 ;
        RECT  9.420 2.075 9.685 2.635 ;
        RECT  9.200 2.075 9.420 2.415 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.755 -0.400 25.080 0.400 ;
        RECT  24.415 -0.400 24.755 0.575 ;
        RECT  23.355 -0.400 24.415 0.400 ;
        RECT  23.015 -0.400 23.355 1.590 ;
        RECT  21.875 -0.400 23.015 0.400 ;
        RECT  21.535 -0.400 21.875 0.575 ;
        RECT  16.815 -0.400 21.535 0.400 ;
        RECT  16.475 -0.400 16.815 0.575 ;
        RECT  15.295 -0.400 16.475 0.400 ;
        RECT  14.955 -0.400 15.295 0.575 ;
        RECT  13.045 -0.400 14.955 0.400 ;
        RECT  12.705 -0.400 13.045 1.270 ;
        RECT  10.385 -0.400 12.705 0.400 ;
        RECT  10.045 -0.400 10.385 0.575 ;
        RECT  6.925 -0.400 10.045 0.400 ;
        RECT  6.585 -0.400 6.925 0.575 ;
        RECT  4.235 -0.400 6.585 0.400 ;
        RECT  3.895 -0.400 4.235 0.575 ;
        RECT  1.120 -0.400 3.895 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.765 4.640 25.080 5.440 ;
        RECT  24.425 4.465 24.765 5.440 ;
        RECT  23.355 4.640 24.425 5.440 ;
        RECT  23.015 3.025 23.355 5.440 ;
        RECT  21.875 4.640 23.015 5.440 ;
        RECT  21.015 4.465 21.875 5.440 ;
        RECT  12.235 4.640 21.015 5.440 ;
        RECT  11.315 4.465 12.235 5.440 ;
        RECT  10.265 4.640 11.315 5.440 ;
        RECT  9.925 4.465 10.265 5.440 ;
        RECT  6.910 4.640 9.925 5.440 ;
        RECT  6.570 4.465 6.910 5.440 ;
        RECT  4.225 4.640 6.570 5.440 ;
        RECT  3.885 4.465 4.225 5.440 ;
        RECT  1.180 4.640 3.885 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.565 2.130 23.505 2.475 ;
        RECT  22.565 1.220 22.635 1.560 ;
        RECT  22.580 3.010 22.635 3.820 ;
        RECT  22.565 3.010 22.580 4.230 ;
        RECT  22.335 1.220 22.565 4.230 ;
        RECT  22.295 1.220 22.335 1.560 ;
        RECT  22.295 3.010 22.335 4.230 ;
        RECT  16.485 4.000 22.295 4.230 ;
        RECT  21.840 2.280 21.970 2.635 ;
        RECT  21.610 0.805 21.840 3.770 ;
        RECT  18.695 0.805 21.610 1.035 ;
        RECT  18.215 3.540 21.610 3.770 ;
        RECT  21.140 1.265 21.370 3.305 ;
        RECT  18.180 1.265 21.140 1.495 ;
        RECT  18.935 3.075 21.140 3.305 ;
        RECT  20.635 1.755 20.865 2.460 ;
        RECT  17.980 2.230 20.635 2.460 ;
        RECT  17.370 1.265 18.180 1.645 ;
        RECT  17.750 2.230 17.980 3.770 ;
        RECT  17.295 0.635 17.945 0.865 ;
        RECT  17.575 2.230 17.750 2.460 ;
        RECT  16.000 3.540 17.750 3.770 ;
        RECT  17.290 2.905 17.520 3.305 ;
        RECT  16.000 1.265 17.370 1.495 ;
        RECT  17.065 0.635 17.295 1.035 ;
        RECT  16.000 3.075 17.290 3.305 ;
        RECT  14.520 0.805 17.065 1.035 ;
        RECT  16.255 4.000 16.485 4.410 ;
        RECT  12.780 4.180 16.255 4.410 ;
        RECT  15.770 1.265 16.000 3.305 ;
        RECT  15.770 3.540 16.000 3.950 ;
        RECT  13.245 3.720 15.770 3.950 ;
        RECT  15.250 2.135 15.480 3.490 ;
        RECT  13.710 3.260 15.250 3.490 ;
        RECT  14.230 2.795 14.575 3.025 ;
        RECT  14.230 0.805 14.520 1.490 ;
        RECT  14.000 0.805 14.230 3.025 ;
        RECT  13.480 1.180 13.710 3.490 ;
        RECT  12.580 2.635 13.480 2.865 ;
        RECT  13.020 1.500 13.250 2.305 ;
        RECT  13.015 3.540 13.245 3.950 ;
        RECT  11.755 1.500 13.020 1.730 ;
        RECT  11.960 3.540 13.015 3.770 ;
        RECT  12.550 4.000 12.780 4.410 ;
        RECT  12.350 2.270 12.580 2.865 ;
        RECT  11.495 4.000 12.550 4.230 ;
        RECT  11.730 3.085 11.960 3.770 ;
        RECT  11.525 1.025 11.755 2.855 ;
        RECT  11.055 3.085 11.730 3.315 ;
        RECT  11.345 1.025 11.525 1.255 ;
        RECT  11.345 2.625 11.525 2.855 ;
        RECT  11.265 3.545 11.495 4.230 ;
        RECT  11.055 1.655 11.275 1.885 ;
        RECT  8.850 3.545 11.265 3.775 ;
        RECT  10.825 1.080 11.055 3.315 ;
        RECT  9.320 4.005 10.895 4.235 ;
        RECT  9.605 1.080 10.825 1.310 ;
        RECT  9.165 3.010 10.825 3.240 ;
        RECT  9.265 0.970 9.605 1.310 ;
        RECT  9.090 4.005 9.320 4.330 ;
        RECT  7.475 4.100 9.090 4.330 ;
        RECT  8.800 1.285 8.850 3.775 ;
        RECT  8.620 1.285 8.800 3.845 ;
        RECT  8.460 3.505 8.620 3.845 ;
        RECT  8.210 1.640 8.330 3.115 ;
        RECT  8.130 1.640 8.210 3.730 ;
        RECT  8.100 1.285 8.130 3.730 ;
        RECT  7.900 1.285 8.100 1.870 ;
        RECT  8.080 2.885 8.100 3.730 ;
        RECT  7.980 2.885 8.080 3.845 ;
        RECT  7.740 3.500 7.980 3.845 ;
        RECT  7.670 2.275 7.865 2.650 ;
        RECT  7.670 0.630 7.805 0.860 ;
        RECT  5.460 3.500 7.740 3.730 ;
        RECT  7.440 0.630 7.670 3.145 ;
        RECT  7.245 4.005 7.475 4.330 ;
        RECT  6.130 0.805 7.440 1.035 ;
        RECT  2.545 4.005 7.245 4.235 ;
        RECT  6.960 1.575 7.190 2.025 ;
        RECT  6.130 1.795 6.960 2.025 ;
        RECT  6.130 2.860 6.295 3.090 ;
        RECT  6.130 1.270 6.265 1.500 ;
        RECT  5.900 0.675 6.130 1.035 ;
        RECT  5.900 1.270 6.130 3.090 ;
        RECT  4.935 0.675 5.900 0.905 ;
        RECT  5.780 2.210 5.900 2.575 ;
        RECT  5.230 1.205 5.460 3.730 ;
        RECT  3.830 3.500 5.230 3.730 ;
        RECT  4.720 1.260 4.950 3.045 ;
        RECT  4.455 1.260 4.720 1.490 ;
        RECT  4.455 2.815 4.720 3.045 ;
        RECT  3.600 0.850 3.830 3.730 ;
        RECT  3.380 0.850 3.600 1.080 ;
        RECT  3.030 3.500 3.600 3.730 ;
        RECT  3.150 0.685 3.380 1.080 ;
        RECT  3.135 1.335 3.365 3.080 ;
        RECT  3.030 0.685 3.150 0.915 ;
        RECT  2.985 1.970 3.135 2.325 ;
        RECT  2.545 1.440 2.665 2.105 ;
        RECT  2.435 1.440 2.545 4.235 ;
        RECT  2.315 1.875 2.435 4.235 ;
        RECT  1.785 3.925 2.015 4.410 ;
        RECT  1.810 1.440 1.920 1.780 ;
        RECT  1.810 3.135 1.840 3.475 ;
        RECT  1.580 1.440 1.810 3.475 ;
        RECT  0.520 3.925 1.785 4.155 ;
        RECT  1.500 3.135 1.580 3.475 ;
        RECT  0.410 1.440 0.520 1.780 ;
        RECT  0.410 3.135 0.520 4.155 ;
        RECT  0.290 1.440 0.410 4.155 ;
        RECT  0.180 1.440 0.290 3.475 ;
    END
END SEDFFHQX4

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFHQXL ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 0.700 1.945 1.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.060 1.105 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.295 1.455 22.300 3.080 ;
        RECT  22.070 1.455 22.295 3.220 ;
        RECT  21.900 1.455 22.070 1.795 ;
        RECT  21.920 2.740 22.070 3.220 ;
        RECT  21.900 2.740 21.920 3.080 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.740 2.305 7.120 2.910 ;
        RECT  6.475 2.330 6.740 2.560 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.485 2.370 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.310 1.770 9.995 2.150 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.560 -0.400 22.440 0.400 ;
        RECT  21.220 -0.400 21.560 0.575 ;
        RECT  20.135 -0.400 21.220 0.400 ;
        RECT  19.795 -0.400 20.135 0.575 ;
        RECT  16.735 -0.400 19.795 0.400 ;
        RECT  16.395 -0.400 16.735 1.720 ;
        RECT  15.295 -0.400 16.395 0.400 ;
        RECT  14.955 -0.400 15.295 1.500 ;
        RECT  13.045 -0.400 14.955 0.400 ;
        RECT  12.705 -0.400 13.045 1.270 ;
        RECT  10.385 -0.400 12.705 0.400 ;
        RECT  10.045 -0.400 10.385 0.575 ;
        RECT  6.925 -0.400 10.045 0.400 ;
        RECT  6.585 -0.400 6.925 0.575 ;
        RECT  4.235 -0.400 6.585 0.400 ;
        RECT  3.895 -0.400 4.235 0.575 ;
        RECT  1.120 -0.400 3.895 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.560 4.640 22.440 5.440 ;
        RECT  21.220 4.465 21.560 5.440 ;
        RECT  20.065 4.640 21.220 5.440 ;
        RECT  19.725 4.465 20.065 5.440 ;
        RECT  12.315 4.640 19.725 5.440 ;
        RECT  11.975 4.465 12.315 5.440 ;
        RECT  10.210 4.640 11.975 5.440 ;
        RECT  9.980 3.725 10.210 5.440 ;
        RECT  6.910 4.640 9.980 5.440 ;
        RECT  6.570 4.465 6.910 5.440 ;
        RECT  4.225 4.640 6.570 5.440 ;
        RECT  3.885 4.465 4.225 5.440 ;
        RECT  1.180 4.640 3.885 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.495 2.100 21.835 2.440 ;
        RECT  20.895 2.210 21.495 2.440 ;
        RECT  20.890 1.225 20.895 1.565 ;
        RECT  20.890 2.210 20.895 3.950 ;
        RECT  20.660 1.225 20.890 3.950 ;
        RECT  20.555 1.225 20.660 1.565 ;
        RECT  20.555 3.140 20.660 3.950 ;
        RECT  19.690 3.590 20.555 3.820 ;
        RECT  20.360 2.280 20.415 2.620 ;
        RECT  20.075 2.280 20.360 2.635 ;
        RECT  19.645 2.405 20.075 2.635 ;
        RECT  19.460 2.870 19.690 3.820 ;
        RECT  19.415 0.895 19.645 2.635 ;
        RECT  19.450 3.590 19.460 3.820 ;
        RECT  19.220 3.590 19.450 4.410 ;
        RECT  19.365 0.895 19.415 1.125 ;
        RECT  19.145 2.405 19.415 2.635 ;
        RECT  19.135 0.730 19.365 1.125 ;
        RECT  12.780 4.180 19.220 4.410 ;
        RECT  18.640 1.385 19.160 1.615 ;
        RECT  18.915 2.405 19.145 3.245 ;
        RECT  18.615 0.730 19.135 0.960 ;
        RECT  18.795 3.015 18.915 3.245 ;
        RECT  18.740 3.015 18.795 3.760 ;
        RECT  18.565 3.015 18.740 3.895 ;
        RECT  18.410 1.385 18.640 2.725 ;
        RECT  18.385 0.630 18.615 0.960 ;
        RECT  18.455 3.420 18.565 3.895 ;
        RECT  17.300 3.665 18.455 3.895 ;
        RECT  17.990 2.495 18.410 2.725 ;
        RECT  17.240 0.630 18.385 0.860 ;
        RECT  17.760 3.095 18.075 3.325 ;
        RECT  17.760 1.095 18.015 1.325 ;
        RECT  17.530 1.095 17.760 3.325 ;
        RECT  15.960 1.975 17.530 2.205 ;
        RECT  17.070 3.085 17.300 3.895 ;
        RECT  16.730 2.495 17.285 2.725 ;
        RECT  17.010 0.630 17.240 1.015 ;
        RECT  16.500 2.495 16.730 3.950 ;
        RECT  13.245 3.720 16.500 3.950 ;
        RECT  15.960 1.160 16.015 1.500 ;
        RECT  15.730 1.160 15.960 3.380 ;
        RECT  15.675 1.160 15.730 1.500 ;
        RECT  15.250 2.135 15.480 3.490 ;
        RECT  13.710 3.260 15.250 3.490 ;
        RECT  14.230 1.215 14.575 1.445 ;
        RECT  14.230 2.795 14.575 3.025 ;
        RECT  14.000 1.215 14.230 3.025 ;
        RECT  13.480 0.970 13.710 3.490 ;
        RECT  12.295 2.325 13.480 2.555 ;
        RECT  13.015 3.540 13.245 3.950 ;
        RECT  13.000 1.500 13.230 1.940 ;
        RECT  11.130 3.540 13.015 3.770 ;
        RECT  11.755 1.500 13.000 1.730 ;
        RECT  12.550 4.005 12.780 4.410 ;
        RECT  10.670 4.005 12.550 4.235 ;
        RECT  11.685 1.125 11.755 2.730 ;
        RECT  11.590 1.070 11.685 2.730 ;
        RECT  11.525 1.070 11.590 3.290 ;
        RECT  11.345 1.070 11.525 1.410 ;
        RECT  11.360 2.500 11.525 3.290 ;
        RECT  10.490 1.655 11.275 1.885 ;
        RECT  10.900 2.795 11.130 3.770 ;
        RECT  10.490 2.795 10.900 3.025 ;
        RECT  10.440 3.260 10.670 4.235 ;
        RECT  10.260 1.080 10.490 3.025 ;
        RECT  8.850 3.260 10.440 3.490 ;
        RECT  9.605 1.080 10.260 1.310 ;
        RECT  9.165 2.795 10.260 3.025 ;
        RECT  9.265 0.970 9.605 1.310 ;
        RECT  7.500 4.125 9.280 4.355 ;
        RECT  8.620 1.285 8.850 3.845 ;
        RECT  8.130 1.640 8.330 3.790 ;
        RECT  8.100 1.285 8.130 3.790 ;
        RECT  7.900 1.285 8.100 1.870 ;
        RECT  7.845 3.500 8.100 3.790 ;
        RECT  7.725 2.275 7.865 2.650 ;
        RECT  5.460 3.500 7.845 3.730 ;
        RECT  7.670 0.630 7.805 0.860 ;
        RECT  7.670 2.275 7.725 3.145 ;
        RECT  7.440 0.630 7.670 3.145 ;
        RECT  7.270 4.005 7.500 4.355 ;
        RECT  6.130 0.805 7.440 1.035 ;
        RECT  7.385 2.805 7.440 3.145 ;
        RECT  2.600 4.005 7.270 4.235 ;
        RECT  6.960 1.575 7.190 2.025 ;
        RECT  6.130 1.795 6.960 2.025 ;
        RECT  6.130 2.805 6.295 3.145 ;
        RECT  6.130 1.270 6.265 1.500 ;
        RECT  5.900 0.675 6.130 1.035 ;
        RECT  5.955 1.270 6.130 3.145 ;
        RECT  5.900 1.270 5.955 3.090 ;
        RECT  4.935 0.675 5.900 0.905 ;
        RECT  5.780 2.210 5.900 2.575 ;
        RECT  5.460 1.205 5.515 1.545 ;
        RECT  5.230 1.205 5.460 3.775 ;
        RECT  5.175 1.205 5.230 1.545 ;
        RECT  3.830 3.545 5.230 3.775 ;
        RECT  4.795 1.260 4.945 3.045 ;
        RECT  4.715 1.205 4.795 3.100 ;
        RECT  4.455 1.205 4.715 1.545 ;
        RECT  4.455 2.760 4.715 3.100 ;
        RECT  3.600 0.850 3.830 3.775 ;
        RECT  3.380 0.850 3.600 1.080 ;
        RECT  3.030 3.545 3.600 3.775 ;
        RECT  3.150 0.685 3.380 1.080 ;
        RECT  3.135 1.335 3.365 3.080 ;
        RECT  3.030 0.685 3.150 0.915 ;
        RECT  2.985 1.970 3.135 2.325 ;
        RECT  2.610 1.440 2.720 1.780 ;
        RECT  2.545 1.440 2.610 2.105 ;
        RECT  2.545 3.445 2.600 4.235 ;
        RECT  2.380 1.440 2.545 4.235 ;
        RECT  2.370 1.875 2.380 4.235 ;
        RECT  2.315 1.875 2.370 3.785 ;
        RECT  2.260 3.445 2.315 3.785 ;
        RECT  2.015 4.070 2.070 4.410 ;
        RECT  1.730 3.925 2.015 4.410 ;
        RECT  1.810 1.440 1.920 1.780 ;
        RECT  1.810 3.135 1.840 3.475 ;
        RECT  1.580 1.440 1.810 3.475 ;
        RECT  0.520 3.925 1.730 4.155 ;
        RECT  1.500 3.135 1.580 3.475 ;
        RECT  0.410 1.440 0.520 1.780 ;
        RECT  0.410 3.135 0.520 4.155 ;
        RECT  0.290 1.440 0.410 4.155 ;
        RECT  0.180 1.440 0.290 3.475 ;
    END
END SEDFFHQX2

MACRO SEDFFHQX1
    CLASS CORE ;
    FOREIGN SEDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFHQXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 0.700 1.945 1.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.060 1.105 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.015 1.360 20.245 3.240 ;
        RECT  19.805 1.360 20.015 1.700 ;
        RECT  19.895 2.900 20.015 3.240 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.740 2.305 7.120 2.910 ;
        RECT  6.475 2.330 6.740 2.560 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.485 2.370 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  9.310 1.770 9.995 2.150 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.585 -0.400 20.460 0.400 ;
        RECT  19.245 -0.400 19.585 0.575 ;
        RECT  18.250 -0.400 19.245 0.400 ;
        RECT  17.910 -0.400 18.250 0.575 ;
        RECT  15.295 -0.400 17.910 0.400 ;
        RECT  14.955 -0.400 15.295 1.615 ;
        RECT  12.965 -0.400 14.955 0.400 ;
        RECT  12.625 -0.400 12.965 1.270 ;
        RECT  10.385 -0.400 12.625 0.400 ;
        RECT  10.045 -0.400 10.385 0.575 ;
        RECT  6.925 -0.400 10.045 0.400 ;
        RECT  6.585 -0.400 6.925 0.575 ;
        RECT  4.235 -0.400 6.585 0.400 ;
        RECT  3.895 -0.400 4.235 0.575 ;
        RECT  1.120 -0.400 3.895 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.680 4.640 20.460 5.440 ;
        RECT  19.250 4.465 19.680 5.440 ;
        RECT  18.210 4.640 19.250 5.440 ;
        RECT  17.870 4.465 18.210 5.440 ;
        RECT  12.315 4.640 17.870 5.440 ;
        RECT  11.975 4.465 12.315 5.440 ;
        RECT  10.210 4.640 11.975 5.440 ;
        RECT  9.980 3.725 10.210 5.440 ;
        RECT  6.910 4.640 9.980 5.440 ;
        RECT  6.570 4.465 6.910 5.440 ;
        RECT  4.225 4.640 6.570 5.440 ;
        RECT  3.885 4.465 4.225 5.440 ;
        RECT  1.180 4.640 3.885 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.415 2.100 19.755 2.440 ;
        RECT  18.920 2.155 19.415 2.385 ;
        RECT  18.920 3.115 18.975 3.925 ;
        RECT  18.885 2.155 18.920 3.925 ;
        RECT  18.655 1.290 18.885 3.925 ;
        RECT  18.545 1.290 18.655 1.630 ;
        RECT  18.635 3.115 18.655 3.925 ;
        RECT  17.835 3.590 18.635 3.820 ;
        RECT  18.025 2.200 18.365 2.540 ;
        RECT  17.730 2.200 18.025 2.430 ;
        RECT  17.835 2.870 17.890 3.210 ;
        RECT  17.605 2.870 17.835 3.820 ;
        RECT  17.670 2.015 17.730 2.430 ;
        RECT  17.440 0.635 17.670 2.430 ;
        RECT  17.550 2.870 17.605 3.210 ;
        RECT  16.880 3.590 17.605 3.820 ;
        RECT  16.680 0.635 17.440 0.865 ;
        RECT  16.915 2.015 17.440 2.245 ;
        RECT  16.980 1.250 17.210 1.625 ;
        RECT  16.440 1.395 16.980 1.625 ;
        RECT  16.880 2.015 16.915 3.240 ;
        RECT  16.685 2.015 16.880 3.360 ;
        RECT  16.650 3.590 16.880 4.410 ;
        RECT  16.650 3.010 16.685 3.360 ;
        RECT  16.450 0.635 16.680 1.125 ;
        RECT  12.780 4.180 16.650 4.410 ;
        RECT  16.420 1.395 16.440 2.810 ;
        RECT  16.210 1.395 16.420 3.950 ;
        RECT  16.190 2.580 16.210 3.950 ;
        RECT  13.245 3.720 16.190 3.950 ;
        RECT  15.730 1.140 15.960 3.275 ;
        RECT  15.250 2.135 15.480 3.490 ;
        RECT  13.710 3.260 15.250 3.490 ;
        RECT  14.245 2.795 14.575 3.025 ;
        RECT  14.245 1.330 14.495 1.560 ;
        RECT  14.015 0.630 14.245 3.025 ;
        RECT  13.480 0.980 13.710 3.490 ;
        RECT  12.295 2.325 13.480 2.555 ;
        RECT  13.015 3.540 13.245 3.950 ;
        RECT  13.000 1.500 13.230 1.940 ;
        RECT  11.130 3.540 13.015 3.770 ;
        RECT  11.755 1.500 13.000 1.730 ;
        RECT  12.550 4.005 12.780 4.410 ;
        RECT  10.670 4.005 12.550 4.235 ;
        RECT  11.590 1.025 11.755 2.730 ;
        RECT  11.525 1.025 11.590 3.290 ;
        RECT  11.265 1.025 11.525 1.255 ;
        RECT  11.360 2.500 11.525 3.290 ;
        RECT  10.455 1.655 11.235 1.885 ;
        RECT  10.900 2.795 11.130 3.770 ;
        RECT  10.455 2.795 10.900 3.025 ;
        RECT  10.440 3.260 10.670 4.235 ;
        RECT  10.225 1.080 10.455 3.025 ;
        RECT  8.850 3.260 10.440 3.490 ;
        RECT  9.605 1.080 10.225 1.310 ;
        RECT  9.165 2.795 10.225 3.025 ;
        RECT  9.265 0.970 9.605 1.310 ;
        RECT  7.500 4.125 9.280 4.355 ;
        RECT  8.620 1.285 8.850 3.845 ;
        RECT  8.130 1.640 8.330 3.790 ;
        RECT  8.100 1.285 8.130 3.790 ;
        RECT  7.900 1.285 8.100 1.870 ;
        RECT  7.845 3.500 8.100 3.790 ;
        RECT  7.670 2.275 7.865 2.650 ;
        RECT  5.460 3.500 7.845 3.730 ;
        RECT  7.670 0.630 7.805 0.860 ;
        RECT  7.440 0.630 7.670 3.145 ;
        RECT  7.270 4.005 7.500 4.355 ;
        RECT  6.130 0.805 7.440 1.035 ;
        RECT  2.545 4.005 7.270 4.235 ;
        RECT  6.960 1.575 7.190 2.025 ;
        RECT  6.130 1.795 6.960 2.025 ;
        RECT  6.130 2.860 6.295 3.090 ;
        RECT  6.130 1.270 6.265 1.500 ;
        RECT  5.900 0.675 6.130 1.035 ;
        RECT  5.900 1.270 6.130 3.090 ;
        RECT  4.935 0.675 5.900 0.905 ;
        RECT  5.780 2.210 5.900 2.575 ;
        RECT  5.230 1.205 5.460 3.730 ;
        RECT  3.830 3.500 5.230 3.730 ;
        RECT  4.720 1.260 4.950 3.045 ;
        RECT  4.455 1.260 4.720 1.490 ;
        RECT  4.455 2.815 4.720 3.045 ;
        RECT  3.600 0.850 3.830 3.730 ;
        RECT  3.380 0.850 3.600 1.080 ;
        RECT  3.030 3.500 3.600 3.730 ;
        RECT  3.150 0.685 3.380 1.080 ;
        RECT  3.135 1.335 3.365 3.080 ;
        RECT  3.030 0.685 3.150 0.915 ;
        RECT  2.985 1.970 3.135 2.325 ;
        RECT  2.545 1.440 2.665 2.105 ;
        RECT  2.435 1.440 2.545 4.235 ;
        RECT  2.315 1.875 2.435 4.235 ;
        RECT  1.785 3.925 2.015 4.410 ;
        RECT  1.810 1.440 1.920 1.780 ;
        RECT  1.810 3.135 1.840 3.475 ;
        RECT  1.580 1.440 1.810 3.475 ;
        RECT  0.520 3.925 1.785 4.155 ;
        RECT  1.500 3.135 1.580 3.475 ;
        RECT  0.410 1.440 0.520 1.780 ;
        RECT  0.410 3.135 0.520 4.155 ;
        RECT  0.290 1.440 0.410 4.155 ;
        RECT  0.180 1.440 0.290 3.475 ;
    END
END SEDFFHQX1

MACRO SDFFTRXL
    CLASS CORE ;
    FOREIGN SDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.420 3.730 2.665 ;
        RECT  2.855 2.405 3.085 2.665 ;
        RECT  2.775 2.420 2.855 2.665 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.925 3.970 3.155 ;
        RECT  2.310 2.925 2.425 3.195 ;
        RECT  2.195 2.335 2.310 3.195 ;
        RECT  2.100 2.335 2.195 3.155 ;
        RECT  2.080 2.200 2.100 3.155 ;
        RECT  1.870 2.200 2.080 2.565 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.820 4.480 2.165 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.150 1.315 14.305 3.160 ;
        RECT  14.080 1.315 14.150 3.270 ;
        RECT  14.075 1.200 14.080 3.270 ;
        RECT  13.785 1.200 14.075 1.545 ;
        RECT  13.810 2.930 14.075 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.555 3.525 13.645 3.755 ;
        RECT  13.325 0.865 13.555 3.970 ;
        RECT  12.605 0.865 13.325 1.095 ;
        RECT  12.890 3.740 13.325 3.970 ;
        RECT  12.550 3.740 12.890 4.080 ;
        RECT  12.375 0.660 12.605 1.095 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.750 1.260 5.180 1.945 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.150 1.180 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.380 -0.400 14.520 0.400 ;
        RECT  13.040 -0.400 13.380 0.575 ;
        RECT  11.900 -0.400 13.040 0.400 ;
        RECT  11.560 -0.400 11.900 0.575 ;
        RECT  9.380 -0.400 11.560 0.400 ;
        RECT  9.040 -0.400 9.380 1.365 ;
        RECT  7.465 -0.400 9.040 0.400 ;
        RECT  7.235 -0.400 7.465 1.060 ;
        RECT  3.410 -0.400 7.235 0.400 ;
        RECT  3.070 -0.400 3.410 0.575 ;
        RECT  1.180 -0.400 3.070 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.590 4.640 14.520 5.440 ;
        RECT  13.535 4.465 13.590 5.440 ;
        RECT  13.305 4.410 13.535 5.440 ;
        RECT  13.250 4.465 13.305 5.440 ;
        RECT  12.130 4.640 13.250 5.440 ;
        RECT  11.790 3.885 12.130 5.440 ;
        RECT  9.850 4.640 11.790 5.440 ;
        RECT  9.510 3.620 9.850 5.440 ;
        RECT  7.390 4.640 9.510 5.440 ;
        RECT  7.335 4.465 7.390 5.440 ;
        RECT  7.105 4.410 7.335 5.440 ;
        RECT  7.050 4.465 7.105 5.440 ;
        RECT  1.210 4.640 7.050 5.440 ;
        RECT  0.790 4.465 1.210 5.440 ;
        RECT  0.000 4.640 0.790 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.890 1.560 13.095 3.020 ;
        RECT  12.865 1.560 12.890 3.130 ;
        RECT  12.700 1.560 12.865 1.790 ;
        RECT  12.550 2.790 12.865 3.130 ;
        RECT  12.360 1.450 12.700 1.790 ;
        RECT  12.320 2.090 12.480 2.430 ;
        RECT  11.750 1.560 12.360 1.790 ;
        RECT  12.140 2.090 12.320 2.690 ;
        RECT  12.090 2.200 12.140 2.690 ;
        RECT  11.075 2.460 12.090 2.690 ;
        RECT  11.520 1.560 11.750 2.230 ;
        RECT  11.410 1.890 11.520 2.230 ;
        RECT  11.075 3.600 11.130 3.940 ;
        RECT  10.845 1.225 11.075 3.940 ;
        RECT  10.615 1.225 10.845 1.455 ;
        RECT  10.790 3.600 10.845 3.940 ;
        RECT  10.385 1.090 10.615 1.455 ;
        RECT  10.155 1.850 10.430 2.190 ;
        RECT  9.925 1.595 10.155 2.975 ;
        RECT  8.670 1.595 9.925 1.825 ;
        RECT  9.255 2.745 9.925 2.975 ;
        RECT  8.210 2.055 9.685 2.395 ;
        RECT  9.025 2.745 9.255 3.190 ;
        RECT  8.445 4.030 8.950 4.260 ;
        RECT  8.440 0.675 8.670 1.825 ;
        RECT  8.215 3.950 8.445 4.260 ;
        RECT  7.710 0.675 8.440 0.905 ;
        RECT  6.605 3.950 8.215 4.180 ;
        RECT  7.990 1.420 8.210 3.135 ;
        RECT  7.980 1.420 7.990 3.190 ;
        RECT  7.870 1.420 7.980 1.760 ;
        RECT  7.650 2.850 7.980 3.190 ;
        RECT  7.560 2.195 7.750 2.540 ;
        RECT  7.065 2.850 7.650 3.080 ;
        RECT  7.520 1.615 7.560 2.540 ;
        RECT  7.330 1.615 7.520 2.425 ;
        RECT  6.265 1.615 7.330 1.845 ;
        RECT  6.835 2.160 7.065 3.080 ;
        RECT  6.305 3.950 6.605 4.410 ;
        RECT  6.255 2.380 6.330 2.720 ;
        RECT  5.705 4.125 6.305 4.410 ;
        RECT  6.255 0.820 6.265 1.845 ;
        RECT  6.160 0.820 6.255 2.720 ;
        RECT  6.025 0.765 6.160 2.720 ;
        RECT  5.820 0.765 6.025 1.105 ;
        RECT  5.990 2.380 6.025 2.720 ;
        RECT  5.705 1.335 5.760 1.675 ;
        RECT  5.475 1.335 5.705 4.410 ;
        RECT  5.420 1.335 5.475 1.675 ;
        RECT  1.685 4.180 5.475 4.410 ;
        RECT  3.875 0.725 5.370 0.955 ;
        RECT  5.045 2.465 5.100 2.805 ;
        RECT  5.045 3.720 5.100 3.950 ;
        RECT  4.815 2.465 5.045 3.950 ;
        RECT  4.760 2.465 4.815 2.805 ;
        RECT  4.705 3.575 4.815 3.950 ;
        RECT  2.345 3.575 4.705 3.805 ;
        RECT  2.870 1.265 4.400 1.495 ;
        RECT  3.645 0.725 3.875 1.035 ;
        RECT  2.545 0.805 3.645 1.035 ;
        RECT  2.640 1.265 2.870 2.000 ;
        RECT  2.530 1.475 2.640 2.000 ;
        RECT  2.315 0.725 2.545 1.035 ;
        RECT  1.920 1.475 2.530 1.705 ;
        RECT  2.005 3.520 2.345 3.860 ;
        RECT  1.710 0.725 2.315 0.955 ;
        RECT  1.640 1.420 1.920 1.760 ;
        RECT  1.640 2.855 1.840 3.085 ;
        RECT  1.455 3.945 1.685 4.410 ;
        RECT  1.580 1.420 1.640 3.085 ;
        RECT  1.410 1.475 1.580 3.085 ;
        RECT  0.520 3.945 1.455 4.175 ;
        RECT  0.415 1.310 0.520 1.650 ;
        RECT  0.415 3.000 0.520 4.175 ;
        RECT  0.290 1.310 0.415 4.175 ;
        RECT  0.185 1.310 0.290 3.340 ;
        RECT  0.180 1.310 0.185 1.650 ;
        RECT  0.180 3.000 0.185 3.340 ;
    END
END SDFFTRXL

MACRO SDFFTRX4
    CLASS CORE ;
    FOREIGN SDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFTRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.600 2.910 4.530 3.200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.235 2.730 5.345 3.070 ;
        RECT  5.005 2.405 5.235 3.070 ;
        RECT  2.210 2.405 5.005 2.635 ;
        RECT  2.120 2.400 2.210 2.635 ;
        RECT  1.870 2.400 2.120 2.740 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.135 2.200 6.190 2.540 ;
        RECT  5.860 2.200 6.135 2.545 ;
        RECT  5.630 1.845 5.860 2.545 ;
        RECT  5.065 1.845 5.630 2.075 ;
        RECT  4.835 1.845 5.065 2.105 ;
        RECT  4.245 1.875 4.835 2.105 ;
        RECT  3.905 1.820 4.245 2.160 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.880 1.260 19.000 2.660 ;
        RECT  18.620 1.260 18.880 3.180 ;
        RECT  18.540 2.840 18.620 3.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.680 1.390 17.700 1.845 ;
        RECT  17.360 1.390 17.680 3.220 ;
        RECT  17.300 1.820 17.360 3.220 ;
        RECT  17.260 2.635 17.300 3.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 1.845 3.085 2.075 ;
        RECT  2.180 1.820 3.080 2.120 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 1.870 1.175 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 -0.400 19.800 0.400 ;
        RECT  19.280 -0.400 19.620 1.000 ;
        RECT  18.340 -0.400 19.280 0.400 ;
        RECT  18.000 -0.400 18.340 1.000 ;
        RECT  17.060 -0.400 18.000 0.400 ;
        RECT  16.720 -0.400 17.060 1.000 ;
        RECT  15.590 -0.400 16.720 0.400 ;
        RECT  15.250 -0.400 15.590 0.575 ;
        RECT  12.900 -0.400 15.250 0.400 ;
        RECT  12.560 -0.400 12.900 1.300 ;
        RECT  10.340 -0.400 12.560 0.400 ;
        RECT  10.000 -0.400 10.340 1.280 ;
        RECT  8.120 -0.400 10.000 0.400 ;
        RECT  7.780 -0.400 8.120 1.410 ;
        RECT  4.680 -0.400 7.780 0.400 ;
        RECT  4.340 -0.400 4.680 0.575 ;
        RECT  1.280 -0.400 4.340 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.520 4.640 19.800 5.440 ;
        RECT  19.180 4.020 19.520 5.440 ;
        RECT  18.240 4.640 19.180 5.440 ;
        RECT  17.900 4.020 18.240 5.440 ;
        RECT  16.960 4.640 17.900 5.440 ;
        RECT  16.620 4.020 16.960 5.440 ;
        RECT  15.620 4.640 16.620 5.440 ;
        RECT  15.280 4.025 15.620 5.440 ;
        RECT  12.940 4.640 15.280 5.440 ;
        RECT  12.600 3.760 12.940 5.440 ;
        RECT  10.340 4.640 12.600 5.440 ;
        RECT  10.000 4.465 10.340 5.440 ;
        RECT  8.660 4.640 10.000 5.440 ;
        RECT  8.605 4.465 8.660 5.440 ;
        RECT  8.375 4.410 8.605 5.440 ;
        RECT  8.320 4.465 8.375 5.440 ;
        RECT  1.280 4.640 8.320 5.440 ;
        RECT  0.940 3.875 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.230 2.210 19.460 3.680 ;
        RECT  16.400 3.450 19.230 3.680 ;
        RECT  16.350 1.395 16.400 3.680 ;
        RECT  16.170 1.290 16.350 3.680 ;
        RECT  16.010 1.290 16.170 1.630 ;
        RECT  15.920 2.940 16.170 3.305 ;
        RECT  15.635 2.010 15.940 2.350 ;
        RECT  15.115 3.075 15.920 3.305 ;
        RECT  15.600 1.350 15.635 2.350 ;
        RECT  15.405 1.350 15.600 2.240 ;
        RECT  14.180 1.350 15.405 1.580 ;
        RECT  14.885 3.075 15.115 3.690 ;
        RECT  14.625 1.820 14.840 2.160 ;
        RECT  14.500 1.820 14.625 4.355 ;
        RECT  14.395 1.875 14.500 4.355 ;
        RECT  13.540 4.125 14.395 4.355 ;
        RECT  14.165 1.240 14.180 1.580 ;
        RECT  13.935 1.240 14.165 3.430 ;
        RECT  13.840 1.240 13.935 1.580 ;
        RECT  11.615 2.095 13.935 2.325 ;
        RECT  13.310 3.215 13.540 4.355 ;
        RECT  12.255 3.215 13.310 3.445 ;
        RECT  12.025 3.215 12.255 4.075 ;
        RECT  9.610 3.845 12.025 4.075 ;
        RECT  11.615 3.275 11.660 3.615 ;
        RECT  11.615 1.025 11.620 1.365 ;
        RECT  11.385 1.025 11.615 3.615 ;
        RECT  11.280 1.025 11.385 1.365 ;
        RECT  11.320 3.275 11.385 3.615 ;
        RECT  10.885 1.595 11.115 2.970 ;
        RECT  9.620 1.595 10.885 1.825 ;
        RECT  9.840 2.740 10.885 2.970 ;
        RECT  9.050 2.115 10.655 2.505 ;
        RECT  9.500 2.735 9.840 3.545 ;
        RECT  9.510 1.105 9.620 1.825 ;
        RECT  9.270 3.790 9.610 4.130 ;
        RECT  9.390 0.630 9.510 1.825 ;
        RECT  9.280 0.630 9.390 1.445 ;
        RECT  8.870 0.630 9.280 0.860 ;
        RECT  8.035 3.900 9.270 4.130 ;
        RECT  8.840 1.340 9.050 2.930 ;
        RECT  8.820 1.230 8.840 2.930 ;
        RECT  8.500 1.230 8.820 1.570 ;
        RECT  8.520 2.700 8.820 2.930 ;
        RECT  8.250 1.910 8.590 2.250 ;
        RECT  8.180 2.700 8.520 3.040 ;
        RECT  7.110 1.965 8.250 2.195 ;
        RECT  7.770 2.735 8.180 2.965 ;
        RECT  7.805 3.900 8.035 4.295 ;
        RECT  6.345 4.065 7.805 4.295 ;
        RECT  7.430 2.700 7.770 3.040 ;
        RECT  6.880 0.845 7.110 3.685 ;
        RECT  6.760 0.845 6.880 1.130 ;
        RECT  6.805 3.455 6.880 3.685 ;
        RECT  6.575 3.455 6.805 3.820 ;
        RECT  6.420 0.790 6.760 1.130 ;
        RECT  6.420 1.360 6.650 3.165 ;
        RECT  6.100 1.360 6.420 1.820 ;
        RECT  6.345 2.935 6.420 3.165 ;
        RECT  6.115 2.935 6.345 4.295 ;
        RECT  2.285 1.360 6.100 1.590 ;
        RECT  5.700 0.790 6.040 1.130 ;
        RECT  5.750 3.820 5.860 4.160 ;
        RECT  5.520 3.455 5.750 4.160 ;
        RECT  2.745 0.845 5.700 1.075 ;
        RECT  2.920 3.455 5.520 3.685 ;
        RECT  4.800 3.960 5.140 4.300 ;
        RECT  2.690 4.015 4.800 4.245 ;
        RECT  2.515 0.685 2.745 1.075 ;
        RECT  2.540 3.310 2.690 4.245 ;
        RECT  2.460 3.255 2.540 4.245 ;
        RECT  2.200 3.255 2.460 3.595 ;
        RECT  2.055 0.865 2.285 1.590 ;
        RECT  2.000 4.065 2.230 4.410 ;
        RECT  0.520 0.865 2.055 1.095 ;
        RECT  1.785 4.065 2.000 4.295 ;
        RECT  1.785 3.020 1.840 3.360 ;
        RECT  1.640 1.420 1.825 1.765 ;
        RECT  1.640 3.020 1.785 4.295 ;
        RECT  1.595 1.420 1.640 4.295 ;
        RECT  1.555 1.535 1.595 4.295 ;
        RECT  1.500 1.535 1.555 3.360 ;
        RECT  1.410 1.535 1.500 3.250 ;
        RECT  0.415 0.845 0.520 1.655 ;
        RECT  0.415 3.050 0.520 3.990 ;
        RECT  0.185 0.845 0.415 3.990 ;
        RECT  0.180 0.845 0.185 1.655 ;
        RECT  0.180 3.050 0.185 3.990 ;
    END
END SDFFTRX4

MACRO SDFFTRX2
    CLASS CORE ;
    FOREIGN SDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFTRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 2.405 3.085 2.635 ;
        RECT  2.790 1.935 3.020 2.635 ;
        RECT  2.780 1.935 2.790 2.380 ;
        RECT  2.680 1.935 2.780 2.165 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.390 1.710 1.840 2.340 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 1.820 3.880 2.370 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.885 1.845 16.945 2.075 ;
        RECT  16.885 3.160 16.890 4.100 ;
        RECT  16.720 1.150 16.885 4.100 ;
        RECT  16.655 1.040 16.720 4.100 ;
        RECT  16.285 1.040 16.655 1.380 ;
        RECT  16.550 3.160 16.655 4.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.185 1.310 15.395 3.130 ;
        RECT  15.165 0.890 15.185 3.130 ;
        RECT  14.845 0.890 15.165 1.540 ;
        RECT  14.735 1.285 14.845 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.600 1.260 5.140 1.675 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.355 1.105 3.195 ;
        RECT  0.645 2.240 0.875 2.585 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.905 -0.400 17.160 0.400 ;
        RECT  15.565 -0.400 15.905 0.950 ;
        RECT  13.765 -0.400 15.565 0.400 ;
        RECT  13.425 -0.400 13.765 1.080 ;
        RECT  11.705 -0.400 13.425 0.400 ;
        RECT  11.365 -0.400 11.705 1.215 ;
        RECT  9.140 -0.400 11.365 0.400 ;
        RECT  8.800 -0.400 9.140 1.270 ;
        RECT  7.225 -0.400 8.800 0.400 ;
        RECT  6.995 -0.400 7.225 0.900 ;
        RECT  3.300 -0.400 6.995 0.400 ;
        RECT  2.960 -0.400 3.300 0.575 ;
        RECT  1.185 -0.400 2.960 0.400 ;
        RECT  0.955 -0.400 1.185 1.450 ;
        RECT  0.000 -0.400 0.955 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.170 4.640 17.160 5.440 ;
        RECT  15.830 4.080 16.170 5.440 ;
        RECT  14.175 4.640 15.830 5.440 ;
        RECT  13.770 4.465 14.175 5.440 ;
        RECT  12.510 4.640 13.770 5.440 ;
        RECT  12.140 4.410 12.510 5.440 ;
        RECT  9.850 4.640 12.140 5.440 ;
        RECT  9.510 4.465 9.850 5.440 ;
        RECT  8.590 4.640 9.510 5.440 ;
        RECT  8.250 4.465 8.590 5.440 ;
        RECT  7.530 4.640 8.250 5.440 ;
        RECT  7.190 4.465 7.530 5.440 ;
        RECT  3.660 4.640 7.190 5.440 ;
        RECT  3.320 4.075 3.660 5.440 ;
        RECT  0.865 4.640 3.320 5.440 ;
        RECT  0.525 4.465 0.865 5.440 ;
        RECT  0.000 4.640 0.525 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.115 2.030 16.330 2.395 ;
        RECT  16.100 2.030 16.115 3.775 ;
        RECT  15.885 2.165 16.100 3.775 ;
        RECT  14.910 3.545 15.885 3.775 ;
        RECT  14.680 1.885 14.910 4.040 ;
        RECT  14.430 1.885 14.680 2.115 ;
        RECT  14.570 3.700 14.680 4.040 ;
        RECT  14.215 2.370 14.445 3.110 ;
        RECT  14.200 0.775 14.430 2.115 ;
        RECT  13.255 2.880 14.215 3.110 ;
        RECT  13.830 1.885 14.200 2.115 ;
        RECT  13.490 1.830 13.830 2.170 ;
        RECT  13.025 1.445 13.255 3.110 ;
        RECT  12.405 1.445 13.025 1.675 ;
        RECT  12.990 2.880 13.025 3.110 ;
        RECT  12.650 2.880 12.990 3.220 ;
        RECT  12.565 1.905 12.795 2.600 ;
        RECT  11.115 2.990 12.650 3.220 ;
        RECT  9.905 1.905 12.565 2.135 ;
        RECT  12.065 0.860 12.405 1.675 ;
        RECT  10.425 1.445 12.065 1.675 ;
        RECT  10.370 2.435 11.165 2.665 ;
        RECT  10.885 2.990 11.115 3.470 ;
        RECT  10.195 0.930 10.425 1.675 ;
        RECT  10.140 2.435 10.370 4.075 ;
        RECT  10.085 0.930 10.195 1.270 ;
        RECT  6.960 3.845 10.140 4.075 ;
        RECT  9.675 1.500 9.905 2.865 ;
        RECT  8.555 1.500 9.675 1.730 ;
        RECT  9.295 2.635 9.675 2.865 ;
        RECT  8.090 1.960 9.445 2.345 ;
        RECT  9.065 2.635 9.295 3.530 ;
        RECT  8.340 0.880 8.555 1.730 ;
        RECT  8.320 0.770 8.340 1.730 ;
        RECT  8.000 0.770 8.320 1.110 ;
        RECT  7.860 1.605 8.090 3.495 ;
        RECT  7.755 0.770 8.000 1.000 ;
        RECT  7.700 1.605 7.860 1.835 ;
        RECT  7.065 3.265 7.860 3.495 ;
        RECT  7.525 0.630 7.755 1.000 ;
        RECT  6.430 2.175 7.630 2.405 ;
        RECT  6.835 2.840 7.065 3.495 ;
        RECT  6.730 3.845 6.960 4.365 ;
        RECT  5.690 4.135 6.730 4.365 ;
        RECT  6.200 0.835 6.430 2.975 ;
        RECT  5.680 0.835 6.200 1.065 ;
        RECT  6.155 2.745 6.200 2.975 ;
        RECT  5.925 2.745 6.155 3.850 ;
        RECT  5.690 1.835 5.970 2.065 ;
        RECT  5.460 1.835 5.690 4.365 ;
        RECT  4.345 4.135 5.460 4.365 ;
        RECT  3.760 0.695 5.220 0.925 ;
        RECT  4.735 2.290 4.965 3.850 ;
        RECT  2.200 3.155 4.735 3.385 ;
        RECT  4.115 3.615 4.345 4.365 ;
        RECT  2.450 1.265 4.260 1.495 ;
        RECT  2.815 3.615 4.115 3.845 ;
        RECT  3.530 0.695 3.760 1.035 ;
        RECT  2.145 0.805 3.530 1.035 ;
        RECT  2.585 3.615 2.815 4.365 ;
        RECT  1.325 4.135 2.585 4.365 ;
        RECT  2.450 2.605 2.550 2.835 ;
        RECT  2.220 1.265 2.450 2.835 ;
        RECT  2.070 1.450 2.220 1.795 ;
        RECT  1.785 2.605 2.220 2.835 ;
        RECT  1.915 0.665 2.145 1.035 ;
        RECT  1.600 0.665 1.915 0.895 ;
        RECT  1.555 2.605 1.785 3.900 ;
        RECT  1.095 3.845 1.325 4.365 ;
        RECT  0.465 3.845 1.095 4.075 ;
        RECT  0.410 1.305 0.520 1.535 ;
        RECT  0.410 3.185 0.465 4.075 ;
        RECT  0.235 1.305 0.410 4.075 ;
        RECT  0.180 1.305 0.235 3.415 ;
    END
END SDFFTRX2

MACRO SDFFTRX1
    CLASS CORE ;
    FOREIGN SDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFTRXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.420 3.730 2.665 ;
        RECT  2.855 2.405 3.085 2.665 ;
        RECT  2.775 2.420 2.855 2.665 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 2.965 3.930 3.195 ;
        RECT  2.120 2.335 2.350 3.195 ;
        RECT  2.100 2.335 2.120 2.565 ;
        RECT  1.870 2.200 2.100 2.565 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.845 4.405 2.165 ;
        RECT  3.590 1.935 4.175 2.165 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.110 1.315 14.305 3.160 ;
        RECT  14.080 1.315 14.110 3.270 ;
        RECT  14.075 1.200 14.080 3.270 ;
        RECT  13.745 1.200 14.075 1.545 ;
        RECT  13.770 2.930 14.075 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.515 3.525 13.645 3.755 ;
        RECT  13.285 0.865 13.515 3.970 ;
        RECT  12.575 0.865 13.285 1.095 ;
        RECT  12.985 3.500 13.285 3.970 ;
        RECT  12.850 3.740 12.985 3.970 ;
        RECT  12.510 3.740 12.850 4.080 ;
        RECT  12.345 0.630 12.575 1.095 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.710 1.260 5.140 1.945 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.150 1.180 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.350 -0.400 14.520 0.400 ;
        RECT  13.010 -0.400 13.350 0.575 ;
        RECT  11.870 -0.400 13.010 0.400 ;
        RECT  11.530 -0.400 11.870 0.575 ;
        RECT  9.350 -0.400 11.530 0.400 ;
        RECT  9.010 -0.400 9.350 1.270 ;
        RECT  7.435 -0.400 9.010 0.400 ;
        RECT  7.205 -0.400 7.435 1.060 ;
        RECT  3.410 -0.400 7.205 0.400 ;
        RECT  3.070 -0.400 3.410 0.575 ;
        RECT  1.180 -0.400 3.070 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.655 4.640 14.520 5.440 ;
        RECT  13.175 4.410 13.655 5.440 ;
        RECT  12.090 4.640 13.175 5.440 ;
        RECT  11.750 4.020 12.090 5.440 ;
        RECT  9.810 4.640 11.750 5.440 ;
        RECT  9.470 3.620 9.810 5.440 ;
        RECT  7.475 4.640 9.470 5.440 ;
        RECT  6.985 4.410 7.475 5.440 ;
        RECT  1.120 4.640 6.985 5.440 ;
        RECT  0.780 4.465 1.120 5.440 ;
        RECT  0.000 4.640 0.780 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.850 1.560 13.055 3.020 ;
        RECT  12.825 1.560 12.850 3.130 ;
        RECT  12.670 1.560 12.825 1.790 ;
        RECT  12.510 2.790 12.825 3.130 ;
        RECT  12.330 1.450 12.670 1.790 ;
        RECT  12.280 2.090 12.440 2.430 ;
        RECT  11.655 1.560 12.330 1.790 ;
        RECT  12.100 2.090 12.280 2.690 ;
        RECT  12.050 2.200 12.100 2.690 ;
        RECT  11.035 2.460 12.050 2.690 ;
        RECT  11.425 1.560 11.655 2.230 ;
        RECT  11.035 3.600 11.090 3.940 ;
        RECT  10.805 1.225 11.035 3.940 ;
        RECT  10.575 1.225 10.805 1.455 ;
        RECT  10.750 3.600 10.805 3.940 ;
        RECT  10.345 1.090 10.575 1.455 ;
        RECT  10.115 1.850 10.380 2.190 ;
        RECT  9.885 1.500 10.115 2.975 ;
        RECT  9.875 1.500 9.885 2.135 ;
        RECT  9.215 2.745 9.885 2.975 ;
        RECT  8.625 1.500 9.875 1.730 ;
        RECT  8.165 1.965 9.645 2.345 ;
        RECT  8.985 2.745 9.215 3.190 ;
        RECT  8.405 4.030 8.910 4.260 ;
        RECT  8.385 0.675 8.625 1.730 ;
        RECT  8.175 3.950 8.405 4.260 ;
        RECT  7.680 0.675 8.385 0.905 ;
        RECT  6.495 3.950 8.175 4.180 ;
        RECT  8.155 1.965 8.165 3.135 ;
        RECT  8.090 1.530 8.155 3.135 ;
        RECT  7.950 1.420 8.090 3.135 ;
        RECT  7.935 1.420 7.950 3.190 ;
        RECT  7.925 1.420 7.935 2.195 ;
        RECT  7.610 2.850 7.935 3.190 ;
        RECT  7.750 1.420 7.925 1.760 ;
        RECT  7.520 2.195 7.695 2.540 ;
        RECT  7.025 2.850 7.610 3.080 ;
        RECT  7.465 1.615 7.520 2.540 ;
        RECT  7.290 1.615 7.465 2.425 ;
        RECT  6.235 1.615 7.290 1.845 ;
        RECT  6.795 2.160 7.025 3.080 ;
        RECT  6.265 3.950 6.495 4.355 ;
        RECT  6.235 2.700 6.290 3.040 ;
        RECT  5.665 4.125 6.265 4.355 ;
        RECT  6.005 0.865 6.235 3.040 ;
        RECT  5.995 0.865 6.005 1.845 ;
        RECT  5.950 2.700 6.005 3.040 ;
        RECT  5.790 0.865 5.995 1.095 ;
        RECT  5.435 1.390 5.665 4.355 ;
        RECT  1.580 4.125 5.435 4.355 ;
        RECT  3.875 0.675 5.330 0.905 ;
        RECT  5.005 2.530 5.060 2.870 ;
        RECT  5.005 3.665 5.060 3.895 ;
        RECT  4.775 2.530 5.005 3.895 ;
        RECT  4.720 2.530 4.775 2.870 ;
        RECT  4.705 3.575 4.775 3.895 ;
        RECT  2.345 3.575 4.705 3.805 ;
        RECT  2.830 1.265 4.360 1.495 ;
        RECT  3.645 0.675 3.875 1.035 ;
        RECT  2.545 0.805 3.645 1.035 ;
        RECT  2.600 1.265 2.830 2.000 ;
        RECT  2.490 1.475 2.600 2.000 ;
        RECT  2.315 0.725 2.545 1.035 ;
        RECT  1.880 1.475 2.490 1.705 ;
        RECT  2.005 3.520 2.345 3.860 ;
        RECT  1.710 0.725 2.315 0.955 ;
        RECT  1.640 1.420 1.880 1.760 ;
        RECT  1.640 2.855 1.840 3.085 ;
        RECT  1.540 1.420 1.640 3.085 ;
        RECT  1.350 3.945 1.580 4.355 ;
        RECT  1.410 1.475 1.540 3.085 ;
        RECT  0.520 3.945 1.350 4.175 ;
        RECT  0.415 1.310 0.520 1.650 ;
        RECT  0.415 2.970 0.520 4.175 ;
        RECT  0.290 1.310 0.415 4.175 ;
        RECT  0.185 1.310 0.290 3.310 ;
        RECT  0.180 1.310 0.185 1.650 ;
        RECT  0.180 2.970 0.185 3.310 ;
    END
END SDFFTRX1

MACRO SDFFSRHQXL
    CLASS CORE ;
    FOREIGN SDFFSRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.680 2.705 18.935 2.935 ;
        RECT  17.500 2.635 17.680 2.965 ;
        RECT  17.270 2.305 17.500 4.045 ;
        RECT  17.265 2.305 17.270 2.935 ;
        RECT  13.925 3.815 17.270 4.045 ;
        RECT  17.095 2.305 17.265 2.535 ;
        RECT  13.885 2.765 13.925 4.045 ;
        RECT  13.775 2.710 13.885 4.045 ;
        RECT  13.695 2.405 13.775 4.045 ;
        RECT  13.545 2.405 13.695 3.240 ;
        RECT  13.415 2.405 13.545 2.635 ;
        RECT  12.965 3.010 13.545 3.240 ;
        RECT  12.735 3.010 12.965 4.405 ;
        RECT  10.275 4.175 12.735 4.405 ;
        RECT  10.045 3.435 10.275 4.405 ;
        RECT  9.350 3.435 10.045 3.665 ;
        RECT  9.120 3.435 9.350 4.410 ;
        RECT  9.025 4.085 9.120 4.410 ;
        RECT  7.445 4.180 9.025 4.410 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.305 2.380 3.820 2.760 ;
        RECT  3.070 2.420 3.305 2.760 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.865 1.285 5.065 1.515 ;
        RECT  4.635 1.285 4.865 2.315 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.725 2.315 16.360 2.855 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.510 1.845 19.585 2.075 ;
        RECT  19.280 1.385 19.510 3.720 ;
        RECT  18.655 1.385 19.280 1.615 ;
        RECT  18.695 3.490 19.280 3.720 ;
        RECT  18.665 3.490 18.695 3.755 ;
        RECT  18.325 3.435 18.665 3.775 ;
        RECT  18.315 1.275 18.655 1.615 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 2.330 2.055 2.765 ;
        RECT  1.455 2.335 1.715 2.765 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.135 1.180 2.575 ;
        RECT  0.645 2.135 1.105 2.635 ;
        RECT  0.640 2.135 0.645 2.575 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.215 -0.400 19.800 0.400 ;
        RECT  16.875 -0.400 17.215 1.615 ;
        RECT  13.455 -0.400 16.875 0.400 ;
        RECT  13.115 -0.400 13.455 0.575 ;
        RECT  10.565 -0.400 13.115 0.400 ;
        RECT  10.225 -0.400 10.565 1.075 ;
        RECT  7.120 -0.400 10.225 0.400 ;
        RECT  6.780 -0.400 7.120 0.900 ;
        RECT  3.475 -0.400 6.780 0.400 ;
        RECT  3.135 -0.400 3.475 0.900 ;
        RECT  1.080 -0.400 3.135 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.455 4.640 19.800 5.440 ;
        RECT  19.115 4.465 19.455 5.440 ;
        RECT  17.325 4.640 19.115 5.440 ;
        RECT  16.985 4.465 17.325 5.440 ;
        RECT  15.800 4.640 16.985 5.440 ;
        RECT  15.460 4.465 15.800 5.440 ;
        RECT  13.465 4.640 15.460 5.440 ;
        RECT  13.235 3.640 13.465 5.440 ;
        RECT  9.810 4.640 13.235 5.440 ;
        RECT  9.580 3.915 9.810 5.440 ;
        RECT  7.115 4.640 9.580 5.440 ;
        RECT  6.775 4.465 7.115 5.440 ;
        RECT  3.040 4.640 6.775 5.440 ;
        RECT  2.810 3.980 3.040 5.440 ;
        RECT  2.700 3.980 2.810 4.210 ;
        RECT  1.595 4.640 2.810 5.440 ;
        RECT  1.175 4.375 1.595 5.440 ;
        RECT  0.000 4.640 1.175 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.080 0.810 19.420 1.150 ;
        RECT  17.935 0.810 19.080 1.040 ;
        RECT  18.840 1.970 18.895 2.310 ;
        RECT  18.555 1.845 18.840 2.310 ;
        RECT  16.860 1.845 18.555 2.075 ;
        RECT  17.705 0.810 17.935 1.555 ;
        RECT  17.595 1.215 17.705 1.555 ;
        RECT  16.630 1.845 16.860 3.525 ;
        RECT  16.345 1.845 16.630 2.075 ;
        RECT  15.340 3.295 16.630 3.525 ;
        RECT  16.115 1.415 16.345 2.075 ;
        RECT  15.610 0.770 15.870 1.000 ;
        RECT  15.380 0.770 15.610 1.135 ;
        RECT  15.340 2.480 15.395 2.820 ;
        RECT  14.880 0.905 15.380 1.135 ;
        RECT  15.110 2.480 15.340 3.525 ;
        RECT  15.055 2.480 15.110 2.820 ;
        RECT  14.730 1.740 15.070 2.080 ;
        RECT  14.650 0.905 14.880 1.505 ;
        RECT  14.385 1.750 14.730 2.015 ;
        RECT  13.920 1.275 14.650 1.505 ;
        RECT  13.955 0.715 14.405 0.945 ;
        RECT  14.155 1.750 14.385 3.580 ;
        RECT  13.100 1.750 14.155 2.015 ;
        RECT  13.725 0.715 13.955 1.035 ;
        RECT  13.365 0.805 13.725 1.035 ;
        RECT  13.135 0.805 13.365 1.280 ;
        RECT  12.500 1.050 13.135 1.280 ;
        RECT  12.760 1.715 13.100 2.055 ;
        RECT  12.270 1.050 12.500 3.255 ;
        RECT  12.100 3.605 12.440 3.945 ;
        RECT  11.785 1.050 12.270 1.280 ;
        RECT  11.675 3.025 12.270 3.255 ;
        RECT  10.735 3.715 12.100 3.945 ;
        RECT  11.805 1.510 12.035 2.795 ;
        RECT  11.365 1.510 11.805 1.740 ;
        RECT  11.195 2.565 11.805 2.795 ;
        RECT  11.285 1.970 11.515 2.310 ;
        RECT  11.135 1.070 11.365 1.740 ;
        RECT  10.735 2.075 11.285 2.310 ;
        RECT  10.965 2.565 11.195 3.480 ;
        RECT  11.025 1.070 11.135 1.410 ;
        RECT  10.505 1.310 10.735 3.945 ;
        RECT  9.765 1.310 10.505 1.540 ;
        RECT  9.530 2.975 10.505 3.205 ;
        RECT  9.920 2.200 10.235 2.540 ;
        RECT  9.895 1.775 9.920 2.540 ;
        RECT  9.690 1.775 9.895 2.485 ;
        RECT  9.605 1.200 9.765 1.540 ;
        RECT  8.460 1.775 9.690 2.005 ;
        RECT  9.425 0.630 9.605 1.540 ;
        RECT  9.375 0.630 9.425 1.485 ;
        RECT  9.070 2.240 9.410 2.580 ;
        RECT  9.265 0.630 9.375 0.970 ;
        RECT  8.885 2.350 9.070 2.580 ;
        RECT  8.655 2.350 8.885 3.845 ;
        RECT  6.295 3.615 8.655 3.845 ;
        RECT  8.425 1.300 8.460 2.005 ;
        RECT  8.195 1.300 8.425 3.270 ;
        RECT  8.120 1.300 8.195 1.640 ;
        RECT  7.775 3.040 8.195 3.270 ;
        RECT  7.735 2.005 7.965 2.380 ;
        RECT  7.435 3.040 7.775 3.380 ;
        RECT  6.080 2.005 7.735 2.235 ;
        RECT  6.820 3.040 7.435 3.270 ;
        RECT  6.590 2.525 6.820 3.270 ;
        RECT  6.385 2.525 6.590 2.755 ;
        RECT  6.065 3.615 6.295 4.345 ;
        RECT  5.885 1.010 6.080 2.735 ;
        RECT  5.325 4.115 6.065 4.345 ;
        RECT  5.850 0.955 5.885 2.735 ;
        RECT  5.545 0.955 5.850 1.295 ;
        RECT  5.785 2.505 5.850 2.735 ;
        RECT  5.555 2.505 5.785 3.825 ;
        RECT  5.325 1.785 5.605 2.125 ;
        RECT  5.265 1.785 5.325 4.345 ;
        RECT  5.095 1.840 5.265 4.345 ;
        RECT  3.500 4.115 5.095 4.345 ;
        RECT  3.935 0.710 4.960 0.940 ;
        RECT  4.525 3.515 4.865 3.855 ;
        RECT  3.960 3.570 4.525 3.800 ;
        RECT  4.400 2.580 4.420 3.125 ;
        RECT  4.400 1.355 4.405 2.100 ;
        RECT  4.190 1.355 4.400 3.125 ;
        RECT  4.175 1.355 4.190 2.810 ;
        RECT  4.170 1.410 4.175 2.810 ;
        RECT  2.735 1.870 4.170 2.100 ;
        RECT  3.730 3.055 3.960 3.800 ;
        RECT  3.705 0.710 3.935 1.640 ;
        RECT  2.100 3.055 3.730 3.285 ;
        RECT  2.100 1.410 3.705 1.640 ;
        RECT  3.270 3.515 3.500 4.345 ;
        RECT  0.520 3.515 3.270 3.745 ;
        RECT  2.395 1.870 2.735 2.660 ;
        RECT  1.860 1.870 2.395 2.100 ;
        RECT  1.630 1.675 1.860 2.100 ;
        RECT  1.140 1.675 1.630 1.905 ;
        RECT  0.460 1.460 0.800 1.800 ;
        RECT  0.410 2.860 0.520 3.745 ;
        RECT  0.410 1.570 0.460 1.800 ;
        RECT  0.290 1.570 0.410 3.745 ;
        RECT  0.180 1.570 0.290 3.200 ;
    END
END SDFFSRHQXL

MACRO SDFFSRHQX4
    CLASS CORE ;
    FOREIGN SDFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRHQXL ;
    SIZE 33.660 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.725 2.495 31.485 2.725 ;
        RECT  26.275 2.085 26.725 2.725 ;
        RECT  26.135 2.495 26.275 2.725 ;
        RECT  25.905 2.495 26.135 4.005 ;
        RECT  21.090 3.775 25.905 4.005 ;
        RECT  21.010 3.315 21.090 4.005 ;
        RECT  21.005 2.370 21.010 4.005 ;
        RECT  20.860 2.315 21.005 4.005 ;
        RECT  20.775 2.315 20.860 3.600 ;
        RECT  20.675 2.405 20.775 2.685 ;
        RECT  20.600 3.195 20.775 3.600 ;
        RECT  20.060 3.370 20.600 3.600 ;
        RECT  19.830 3.370 20.060 4.155 ;
        RECT  12.480 3.925 19.830 4.155 ;
        RECT  12.250 3.580 12.480 4.155 ;
        RECT  11.095 3.580 12.250 3.810 ;
        RECT  10.865 3.580 11.095 4.015 ;
        RECT  8.630 3.785 10.865 4.015 ;
        RECT  8.400 3.785 8.630 4.155 ;
        RECT  8.090 3.925 8.400 4.155 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.825 1.815 3.830 2.045 ;
        RECT  3.165 1.695 3.825 2.125 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.760 5.085 1.990 ;
        RECT  4.175 1.760 4.405 2.075 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.545 2.315 24.235 2.545 ;
        RECT  23.315 2.315 23.545 2.635 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  33.520 3.025 33.525 3.835 ;
        RECT  33.515 2.380 33.520 3.835 ;
        RECT  33.140 1.370 33.515 3.835 ;
        RECT  32.760 1.370 33.140 1.600 ;
        RECT  32.450 3.025 33.140 3.835 ;
        RECT  32.125 1.260 32.760 1.600 ;
        RECT  31.350 3.025 32.450 3.375 ;
        RECT  31.320 1.315 32.125 1.600 ;
        RECT  31.010 3.025 31.350 3.835 ;
        RECT  30.980 1.260 31.320 1.600 ;
        RECT  29.560 3.025 31.010 3.375 ;
        RECT  30.805 1.260 30.980 1.545 ;
        RECT  29.915 1.315 30.805 1.545 ;
        RECT  29.880 1.260 29.915 1.545 ;
        RECT  29.540 1.260 29.880 1.600 ;
        RECT  29.350 3.025 29.560 3.525 ;
        RECT  29.010 3.025 29.350 3.880 ;
        RECT  26.920 3.025 29.010 3.375 ;
        RECT  26.710 3.025 26.920 3.525 ;
        RECT  26.370 3.025 26.710 3.880 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 1.775 2.635 2.635 ;
        RECT  1.540 2.405 2.405 2.635 ;
        RECT  1.300 2.195 1.540 2.635 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.880 0.520 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  28.460 -0.400 33.660 0.400 ;
        RECT  28.120 -0.400 28.460 0.895 ;
        RECT  26.975 -0.400 28.120 0.400 ;
        RECT  26.635 -0.400 26.975 0.895 ;
        RECT  25.400 -0.400 26.635 0.400 ;
        RECT  25.060 -0.400 25.400 1.355 ;
        RECT  23.880 -0.400 25.060 0.400 ;
        RECT  23.540 -0.400 23.880 1.795 ;
        RECT  20.775 -0.400 23.540 0.400 ;
        RECT  20.435 -0.400 20.775 0.575 ;
        RECT  15.590 -0.400 20.435 0.400 ;
        RECT  15.250 -0.400 15.590 0.815 ;
        RECT  14.055 -0.400 15.250 0.400 ;
        RECT  13.715 -0.400 14.055 0.815 ;
        RECT  13.130 -0.400 13.715 0.400 ;
        RECT  12.790 -0.400 13.130 1.090 ;
        RECT  7.805 -0.400 12.790 0.400 ;
        RECT  7.465 -0.400 7.805 0.870 ;
        RECT  4.045 -0.400 7.465 0.400 ;
        RECT  3.815 -0.400 4.045 0.870 ;
        RECT  1.580 -0.400 3.815 0.400 ;
        RECT  1.240 -0.400 1.580 0.575 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  32.070 4.640 33.660 5.440 ;
        RECT  31.730 3.665 32.070 5.440 ;
        RECT  30.630 4.640 31.730 5.440 ;
        RECT  30.290 3.670 30.630 5.440 ;
        RECT  28.030 4.640 30.290 5.440 ;
        RECT  27.690 3.740 28.030 5.440 ;
        RECT  25.070 4.640 27.690 5.440 ;
        RECT  24.730 4.465 25.070 5.440 ;
        RECT  23.485 4.640 24.730 5.440 ;
        RECT  23.145 4.465 23.485 5.440 ;
        RECT  20.625 4.640 23.145 5.440 ;
        RECT  20.395 3.830 20.625 5.440 ;
        RECT  11.665 4.640 20.395 5.440 ;
        RECT  11.325 4.090 11.665 5.440 ;
        RECT  9.335 4.640 11.325 5.440 ;
        RECT  8.995 4.465 9.335 5.440 ;
        RECT  7.840 4.640 8.995 5.440 ;
        RECT  7.610 3.755 7.840 5.440 ;
        RECT  3.115 4.640 7.610 5.440 ;
        RECT  2.775 4.015 3.115 5.440 ;
        RECT  0.520 4.640 2.775 5.440 ;
        RECT  0.180 2.980 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  33.140 0.710 33.480 1.050 ;
        RECT  32.040 0.765 33.140 0.995 ;
        RECT  31.815 1.960 32.625 2.300 ;
        RECT  31.700 0.690 32.040 1.030 ;
        RECT  27.280 2.015 31.815 2.245 ;
        RECT  30.600 0.745 31.700 0.975 ;
        RECT  30.260 0.690 30.600 1.030 ;
        RECT  29.160 0.745 30.260 0.975 ;
        RECT  28.930 0.745 29.160 1.355 ;
        RECT  28.820 1.015 28.930 1.355 ;
        RECT  27.735 1.125 28.820 1.355 ;
        RECT  27.395 0.945 27.735 1.355 ;
        RECT  26.255 1.125 27.395 1.355 ;
        RECT  27.050 1.585 27.280 2.245 ;
        RECT  25.670 1.585 27.050 1.815 ;
        RECT  25.915 1.015 26.255 1.355 ;
        RECT  25.515 1.585 25.670 2.590 ;
        RECT  25.440 1.585 25.515 2.645 ;
        RECT  25.175 2.305 25.440 2.645 ;
        RECT  24.705 2.360 25.175 2.590 ;
        RECT  24.700 1.275 24.705 2.590 ;
        RECT  24.600 1.275 24.700 3.420 ;
        RECT  24.470 0.985 24.600 3.420 ;
        RECT  24.260 0.985 24.470 1.795 ;
        RECT  24.270 3.190 24.470 3.420 ;
        RECT  23.930 3.190 24.270 3.530 ;
        RECT  22.835 3.245 23.930 3.475 ;
        RECT  22.895 0.750 23.125 1.425 ;
        RECT  21.795 0.750 22.895 0.980 ;
        RECT  22.605 2.180 22.835 3.475 ;
        RECT  22.145 1.215 22.375 2.655 ;
        RECT  22.035 1.215 22.145 1.620 ;
        RECT  21.550 2.425 22.145 2.655 ;
        RECT  20.305 1.390 22.035 1.620 ;
        RECT  19.675 1.850 21.885 2.080 ;
        RECT  21.565 0.750 21.795 1.155 ;
        RECT  21.235 0.925 21.565 1.155 ;
        RECT  21.320 2.425 21.550 3.190 ;
        RECT  20.075 1.215 20.305 1.620 ;
        RECT  19.445 0.715 19.675 3.135 ;
        RECT  12.990 3.445 19.475 3.675 ;
        RECT  19.060 0.715 19.445 1.025 ;
        RECT  16.590 2.905 19.445 3.135 ;
        RECT  18.550 0.795 19.060 1.025 ;
        RECT  18.320 0.795 18.550 1.585 ;
        RECT  17.245 0.795 18.320 1.025 ;
        RECT  17.595 1.460 17.825 2.085 ;
        RECT  16.420 1.855 17.595 2.085 ;
        RECT  17.015 0.795 17.245 1.590 ;
        RECT  16.815 1.360 17.015 1.590 ;
        RECT  16.050 0.735 16.720 0.965 ;
        RECT  16.245 1.515 16.420 2.085 ;
        RECT  16.015 1.515 16.245 3.135 ;
        RECT  15.820 0.735 16.050 1.280 ;
        RECT  14.475 1.515 16.015 1.745 ;
        RECT  13.220 2.905 16.015 3.135 ;
        RECT  14.190 1.050 15.820 1.280 ;
        RECT  13.960 1.050 14.190 2.650 ;
        RECT  12.100 1.385 13.960 1.615 ;
        RECT  12.990 2.420 13.960 2.650 ;
        RECT  12.525 1.925 13.515 2.155 ;
        RECT  12.760 2.420 12.990 3.675 ;
        RECT  11.945 3.120 12.760 3.350 ;
        RECT  12.295 1.925 12.525 2.735 ;
        RECT  10.635 2.505 12.295 2.735 ;
        RECT  11.870 0.635 12.100 1.615 ;
        RECT  11.095 2.025 12.065 2.255 ;
        RECT  11.330 0.635 11.560 1.280 ;
        RECT  9.715 0.635 11.330 0.865 ;
        RECT  10.865 1.100 11.095 2.255 ;
        RECT  10.175 1.100 10.865 1.330 ;
        RECT  10.405 1.560 10.635 3.525 ;
        RECT  7.505 3.295 10.405 3.525 ;
        RECT  9.945 1.100 10.175 3.005 ;
        RECT  8.065 2.775 9.945 3.005 ;
        RECT  9.485 0.635 9.715 1.835 ;
        RECT  8.370 1.315 9.485 1.545 ;
        RECT  8.980 2.250 9.285 2.480 ;
        RECT  8.750 1.935 8.980 2.480 ;
        RECT  7.580 1.935 8.750 2.165 ;
        RECT  8.030 1.315 8.370 1.655 ;
        RECT  7.835 2.400 8.065 3.005 ;
        RECT  6.935 2.400 7.835 2.630 ;
        RECT  7.350 1.345 7.580 2.165 ;
        RECT  7.275 2.860 7.505 3.525 ;
        RECT  6.475 1.345 7.350 1.575 ;
        RECT  7.165 2.860 7.275 3.200 ;
        RECT  6.705 2.400 6.935 4.230 ;
        RECT  6.010 4.000 6.705 4.230 ;
        RECT  6.445 1.345 6.475 3.695 ;
        RECT  6.245 0.925 6.445 3.695 ;
        RECT  6.215 0.925 6.245 1.575 ;
        RECT  6.105 0.925 6.215 1.265 ;
        RECT  5.780 1.830 6.010 4.230 ;
        RECT  3.585 4.000 5.780 4.230 ;
        RECT  4.505 0.710 5.720 0.940 ;
        RECT  4.215 3.465 5.550 3.695 ;
        RECT  5.315 1.295 5.545 2.975 ;
        RECT  4.965 1.295 5.315 1.525 ;
        RECT  4.705 2.745 5.315 2.975 ;
        RECT  4.735 1.170 4.965 1.525 ;
        RECT  4.475 2.490 4.705 2.975 ;
        RECT  4.275 0.710 4.505 1.385 ;
        RECT  3.080 2.490 4.475 2.720 ;
        RECT  2.930 1.155 4.275 1.385 ;
        RECT  3.985 3.025 4.215 3.695 ;
        RECT  1.790 3.025 3.985 3.255 ;
        RECT  3.355 3.555 3.585 4.230 ;
        RECT  2.530 3.555 3.355 3.785 ;
        RECT  2.590 1.100 2.930 1.440 ;
        RECT  2.300 3.555 2.530 4.190 ;
        RECT  1.240 3.960 2.300 4.190 ;
        RECT  1.505 3.025 1.790 3.550 ;
        RECT  1.450 3.210 1.505 3.550 ;
        RECT  0.980 3.960 1.240 4.300 ;
        RECT  0.900 1.280 0.980 4.300 ;
        RECT  0.750 1.280 0.900 4.245 ;
        RECT  0.620 1.280 0.750 1.510 ;
        RECT  0.280 0.690 0.620 1.510 ;
    END
END SDFFSRHQX4

MACRO SDFFSRHQX2
    CLASS CORE ;
    FOREIGN SDFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRHQXL ;
    SIZE 25.080 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.245 2.495 22.575 2.725 ;
        RECT  20.015 2.405 20.245 2.725 ;
        RECT  19.765 2.410 20.015 2.725 ;
        RECT  19.535 2.410 19.765 4.005 ;
        RECT  19.510 2.410 19.535 2.640 ;
        RECT  19.355 3.755 19.535 4.005 ;
        RECT  16.210 3.775 19.355 4.005 ;
        RECT  16.210 2.610 16.370 2.840 ;
        RECT  15.980 2.610 16.210 4.005 ;
        RECT  15.155 2.610 15.980 2.840 ;
        RECT  14.925 2.610 15.155 4.315 ;
        RECT  14.735 3.955 14.925 4.315 ;
        RECT  10.260 3.955 14.735 4.185 ;
        RECT  10.030 3.500 10.260 4.185 ;
        RECT  9.340 3.500 10.030 3.730 ;
        RECT  9.110 3.500 9.340 4.290 ;
        RECT  7.325 4.060 9.110 4.290 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 1.750 3.860 2.135 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.685 2.965 1.765 3.195 ;
        RECT  1.235 2.460 1.685 3.220 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.270 1.725 18.310 2.695 ;
        RECT  17.990 1.685 18.270 2.695 ;
        RECT  17.930 1.685 17.990 2.025 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.205 1.370 24.210 3.195 ;
        RECT  23.980 1.370 24.205 3.205 ;
        RECT  23.915 1.370 23.980 1.600 ;
        RECT  23.975 2.965 23.980 3.205 ;
        RECT  22.840 2.975 23.975 3.205 ;
        RECT  23.575 1.260 23.915 1.600 ;
        RECT  23.545 1.285 23.575 1.600 ;
        RECT  22.655 1.370 23.545 1.600 ;
        RECT  22.500 2.975 22.840 3.905 ;
        RECT  22.045 1.260 22.655 1.600 ;
        RECT  20.770 2.975 22.500 3.205 ;
        RECT  20.485 2.975 20.770 4.010 ;
        RECT  20.430 3.190 20.485 4.010 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 2.300 2.495 2.725 ;
        RECT  1.920 2.365 1.925 2.705 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.850 0.520 2.730 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.905 -0.400 25.080 0.400 ;
        RECT  20.565 -0.400 20.905 1.220 ;
        RECT  18.840 -0.400 20.565 0.400 ;
        RECT  18.500 -0.400 18.840 1.455 ;
        RECT  15.815 -0.400 18.500 0.400 ;
        RECT  15.475 -0.400 15.815 0.575 ;
        RECT  11.840 -0.400 15.475 0.400 ;
        RECT  11.500 -0.400 11.840 0.815 ;
        RECT  10.370 -0.400 11.500 0.400 ;
        RECT  10.030 -0.400 10.370 0.820 ;
        RECT  6.985 -0.400 10.030 0.400 ;
        RECT  6.645 -0.400 6.985 1.595 ;
        RECT  3.540 -0.400 6.645 0.400 ;
        RECT  3.200 -0.400 3.540 0.870 ;
        RECT  1.340 -0.400 3.200 0.400 ;
        RECT  1.000 -0.400 1.340 0.575 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.560 4.640 25.080 5.440 ;
        RECT  23.220 3.530 23.560 5.440 ;
        RECT  22.120 4.640 23.220 5.440 ;
        RECT  21.780 3.530 22.120 5.440 ;
        RECT  19.400 4.640 21.780 5.440 ;
        RECT  19.060 4.465 19.400 5.440 ;
        RECT  17.990 4.640 19.060 5.440 ;
        RECT  17.650 4.465 17.990 5.440 ;
        RECT  15.745 4.640 17.650 5.440 ;
        RECT  15.515 3.600 15.745 5.440 ;
        RECT  9.800 4.640 15.515 5.440 ;
        RECT  9.570 3.960 9.800 5.440 ;
        RECT  7.065 4.640 9.570 5.440 ;
        RECT  6.835 3.960 7.065 5.440 ;
        RECT  3.335 4.640 6.835 5.440 ;
        RECT  2.995 3.910 3.335 5.440 ;
        RECT  1.285 4.640 2.995 5.440 ;
        RECT  1.055 3.910 1.285 5.440 ;
        RECT  0.905 3.910 1.055 4.140 ;
        RECT  0.000 4.640 1.055 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  24.675 1.125 24.785 1.465 ;
        RECT  24.445 0.800 24.675 1.465 ;
        RECT  23.150 0.800 24.445 1.030 ;
        RECT  23.515 1.915 23.745 2.350 ;
        RECT  19.565 1.915 23.515 2.145 ;
        RECT  22.810 0.690 23.150 1.030 ;
        RECT  21.665 0.800 22.810 1.030 ;
        RECT  21.610 0.800 21.665 1.490 ;
        RECT  21.435 0.800 21.610 1.685 ;
        RECT  21.325 1.150 21.435 1.685 ;
        RECT  20.105 1.455 21.325 1.685 ;
        RECT  19.875 0.750 20.105 1.685 ;
        RECT  19.765 0.750 19.875 1.090 ;
        RECT  19.225 1.460 19.565 2.145 ;
        RECT  19.105 1.915 19.225 2.145 ;
        RECT  19.105 2.415 19.160 2.755 ;
        RECT  19.050 1.915 19.105 2.755 ;
        RECT  18.875 1.915 19.050 3.155 ;
        RECT  18.820 2.415 18.875 3.155 ;
        RECT  18.750 2.925 18.820 3.155 ;
        RECT  18.465 2.925 18.750 3.450 ;
        RECT  18.410 3.110 18.465 3.450 ;
        RECT  17.745 3.165 18.410 3.395 ;
        RECT  17.890 1.150 18.140 1.380 ;
        RECT  17.660 0.825 17.890 1.380 ;
        RECT  17.515 2.420 17.745 3.395 ;
        RECT  16.180 0.825 17.660 1.055 ;
        RECT  17.335 2.420 17.515 2.650 ;
        RECT  17.265 1.345 17.320 1.575 ;
        RECT  17.075 1.285 17.265 1.575 ;
        RECT  16.845 1.285 17.075 3.300 ;
        RECT  15.495 1.285 16.845 1.515 ;
        RECT  16.670 3.070 16.845 3.300 ;
        RECT  16.440 3.070 16.670 3.460 ;
        RECT  16.385 1.850 16.615 2.325 ;
        RECT  14.390 2.095 16.385 2.325 ;
        RECT  15.265 1.285 15.495 1.805 ;
        RECT  15.060 1.575 15.265 1.805 ;
        RECT  14.020 3.330 14.690 3.560 ;
        RECT  14.315 2.795 14.635 3.025 ;
        RECT  14.390 0.690 14.445 0.920 ;
        RECT  14.315 0.690 14.390 2.325 ;
        RECT  14.085 0.690 14.315 3.025 ;
        RECT  13.285 0.795 14.085 1.025 ;
        RECT  13.350 2.795 14.085 3.025 ;
        RECT  13.790 3.330 14.020 3.645 ;
        RECT  13.620 1.460 13.850 2.045 ;
        RECT  10.720 3.415 13.790 3.645 ;
        RECT  12.500 1.815 13.620 2.045 ;
        RECT  13.010 2.740 13.350 3.080 ;
        RECT  13.055 0.795 13.285 1.585 ;
        RECT  12.835 1.355 13.055 1.585 ;
        RECT  12.430 0.750 12.725 0.980 ;
        RECT  12.240 2.740 12.580 3.080 ;
        RECT  12.110 1.515 12.500 2.045 ;
        RECT  12.200 0.750 12.430 1.280 ;
        RECT  11.180 2.795 12.240 3.025 ;
        RECT  10.505 1.050 12.200 1.280 ;
        RECT  11.180 1.815 12.110 2.045 ;
        RECT  10.950 1.515 11.180 3.080 ;
        RECT  10.735 1.515 10.950 1.745 ;
        RECT  10.505 3.015 10.720 3.645 ;
        RECT  10.490 1.050 10.505 3.645 ;
        RECT  10.275 1.050 10.490 3.245 ;
        RECT  9.570 1.255 10.275 1.485 ;
        RECT  9.580 3.015 10.275 3.245 ;
        RECT  9.815 1.770 10.045 2.520 ;
        RECT  8.415 1.770 9.815 2.000 ;
        RECT  9.460 1.200 9.570 1.540 ;
        RECT  9.230 0.655 9.460 1.540 ;
        RECT  8.875 2.235 9.395 2.465 ;
        RECT  9.060 0.655 9.230 0.885 ;
        RECT  8.645 2.235 8.875 3.675 ;
        RECT  6.110 3.445 8.645 3.675 ;
        RECT  8.305 1.445 8.415 3.215 ;
        RECT  8.185 1.390 8.305 3.215 ;
        RECT  7.965 1.390 8.185 1.730 ;
        RECT  7.055 2.985 8.185 3.215 ;
        RECT  5.655 2.115 7.950 2.345 ;
        RECT  6.825 2.595 7.055 3.215 ;
        RECT  6.500 2.595 6.825 2.825 ;
        RECT  5.880 3.030 6.110 4.410 ;
        RECT  5.180 4.180 5.880 4.410 ;
        RECT  5.645 0.745 5.655 2.345 ;
        RECT  5.415 0.745 5.645 3.910 ;
        RECT  5.280 0.745 5.415 0.975 ;
        RECT  4.950 1.985 5.180 4.410 ;
        RECT  4.760 1.985 4.950 2.215 ;
        RECT  3.800 4.180 4.950 4.410 ;
        RECT  4.005 0.690 4.815 0.920 ;
        RECT  4.490 2.495 4.720 3.030 ;
        RECT  4.380 3.475 4.720 3.815 ;
        RECT  4.465 1.425 4.645 1.655 ;
        RECT  4.465 2.495 4.490 2.735 ;
        RECT  4.235 1.425 4.465 2.735 ;
        RECT  4.260 3.475 4.380 3.705 ;
        RECT  4.030 2.975 4.260 3.705 ;
        RECT  2.960 2.505 4.235 2.735 ;
        RECT  2.270 2.975 4.030 3.205 ;
        RECT  3.775 0.690 4.005 1.500 ;
        RECT  3.570 3.450 3.800 4.410 ;
        RECT  2.540 1.270 3.775 1.500 ;
        RECT  0.980 3.450 3.570 3.680 ;
        RECT  2.730 1.815 2.960 2.735 ;
        RECT  1.250 1.815 2.730 2.045 ;
        RECT  2.200 1.215 2.540 1.555 ;
        RECT  0.750 1.145 0.980 3.680 ;
        RECT  0.520 1.145 0.750 1.375 ;
        RECT  0.520 3.330 0.750 3.680 ;
        RECT  0.180 1.035 0.520 1.375 ;
        RECT  0.180 3.330 0.520 4.150 ;
    END
END SDFFSRHQX2

MACRO SDFFSRHQX1
    CLASS CORE ;
    FOREIGN SDFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRHQXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.680 2.705 18.935 2.935 ;
        RECT  17.500 2.705 17.680 2.965 ;
        RECT  17.270 2.305 17.500 4.045 ;
        RECT  17.265 2.305 17.270 2.935 ;
        RECT  13.925 3.815 17.270 4.045 ;
        RECT  17.095 2.305 17.265 2.535 ;
        RECT  13.885 2.765 13.925 4.045 ;
        RECT  13.775 2.710 13.885 4.045 ;
        RECT  13.695 2.405 13.775 4.045 ;
        RECT  13.545 2.405 13.695 3.240 ;
        RECT  13.415 2.405 13.545 2.635 ;
        RECT  12.965 3.010 13.545 3.240 ;
        RECT  12.735 3.010 12.965 4.365 ;
        RECT  10.275 4.135 12.735 4.365 ;
        RECT  10.045 3.445 10.275 4.365 ;
        RECT  9.350 3.445 10.045 3.675 ;
        RECT  9.120 3.445 9.350 4.410 ;
        RECT  9.025 4.085 9.120 4.410 ;
        RECT  7.445 4.180 9.025 4.410 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.305 2.380 3.820 2.760 ;
        RECT  3.070 2.420 3.305 2.760 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.875 1.285 5.065 1.515 ;
        RECT  4.645 1.285 4.875 2.315 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.065 2.405 16.285 2.635 ;
        RECT  15.835 2.405 16.065 3.020 ;
        RECT  15.725 2.680 15.835 3.020 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.510 1.845 19.585 2.075 ;
        RECT  19.280 1.510 19.510 3.460 ;
        RECT  18.570 1.510 19.280 1.740 ;
        RECT  18.665 3.230 19.280 3.460 ;
        RECT  18.325 3.230 18.665 4.040 ;
        RECT  18.285 1.275 18.570 1.740 ;
        RECT  18.230 1.275 18.285 1.615 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 2.350 2.055 2.790 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.845 1.105 2.540 ;
        RECT  0.645 2.050 0.875 2.540 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.130 -0.400 19.800 0.400 ;
        RECT  16.790 -0.400 17.130 1.615 ;
        RECT  13.455 -0.400 16.790 0.400 ;
        RECT  13.115 -0.400 13.455 0.575 ;
        RECT  10.565 -0.400 13.115 0.400 ;
        RECT  10.225 -0.400 10.565 1.075 ;
        RECT  7.120 -0.400 10.225 0.400 ;
        RECT  6.780 -0.400 7.120 0.900 ;
        RECT  3.390 -0.400 6.780 0.400 ;
        RECT  3.050 -0.400 3.390 0.900 ;
        RECT  1.080 -0.400 3.050 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.455 4.640 19.800 5.440 ;
        RECT  19.115 4.465 19.455 5.440 ;
        RECT  17.325 4.640 19.115 5.440 ;
        RECT  16.985 4.465 17.325 5.440 ;
        RECT  15.600 4.640 16.985 5.440 ;
        RECT  15.260 4.465 15.600 5.440 ;
        RECT  13.465 4.640 15.260 5.440 ;
        RECT  13.235 3.640 13.465 5.440 ;
        RECT  9.810 4.640 13.235 5.440 ;
        RECT  9.580 3.915 9.810 5.440 ;
        RECT  7.115 4.640 9.580 5.440 ;
        RECT  6.775 4.465 7.115 5.440 ;
        RECT  3.040 4.640 6.775 5.440 ;
        RECT  2.810 3.980 3.040 5.440 ;
        RECT  2.700 3.980 2.810 4.210 ;
        RECT  1.595 4.640 2.810 5.440 ;
        RECT  1.175 4.375 1.595 5.440 ;
        RECT  0.000 4.640 1.175 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.280 0.940 19.335 1.280 ;
        RECT  18.995 0.810 19.280 1.280 ;
        RECT  17.850 0.810 18.995 1.040 ;
        RECT  18.555 1.970 18.895 2.310 ;
        RECT  17.990 1.970 18.555 2.205 ;
        RECT  17.730 1.845 17.990 2.205 ;
        RECT  17.620 0.810 17.850 1.375 ;
        RECT  16.860 1.845 17.730 2.075 ;
        RECT  17.510 1.035 17.620 1.375 ;
        RECT  16.860 2.920 16.915 3.260 ;
        RECT  16.805 1.845 16.860 3.260 ;
        RECT  16.630 1.845 16.805 3.525 ;
        RECT  16.370 1.845 16.630 2.075 ;
        RECT  16.575 2.920 16.630 3.525 ;
        RECT  15.340 3.295 16.575 3.525 ;
        RECT  16.140 1.415 16.370 2.075 ;
        RECT  16.030 1.415 16.140 1.755 ;
        RECT  15.610 0.770 15.870 1.000 ;
        RECT  15.380 0.770 15.610 1.135 ;
        RECT  15.340 2.670 15.395 3.010 ;
        RECT  14.880 0.905 15.380 1.135 ;
        RECT  15.110 2.670 15.340 3.525 ;
        RECT  15.055 2.670 15.110 3.010 ;
        RECT  14.730 1.740 15.070 2.080 ;
        RECT  14.650 0.905 14.880 1.505 ;
        RECT  14.385 1.750 14.730 2.015 ;
        RECT  13.920 1.275 14.650 1.505 ;
        RECT  13.955 0.730 14.405 0.960 ;
        RECT  14.155 1.750 14.385 3.580 ;
        RECT  13.070 1.750 14.155 2.015 ;
        RECT  13.725 0.730 13.955 1.035 ;
        RECT  13.365 0.805 13.725 1.035 ;
        RECT  13.135 0.805 13.365 1.185 ;
        RECT  12.495 0.955 13.135 1.185 ;
        RECT  12.730 1.715 13.070 2.055 ;
        RECT  12.265 0.955 12.495 3.225 ;
        RECT  10.735 3.615 12.440 3.845 ;
        RECT  11.745 0.955 12.265 1.185 ;
        RECT  11.760 2.995 12.265 3.225 ;
        RECT  11.805 1.415 12.035 2.710 ;
        RECT  11.325 1.415 11.805 1.645 ;
        RECT  11.195 2.480 11.805 2.710 ;
        RECT  11.230 1.905 11.570 2.245 ;
        RECT  11.040 1.280 11.325 1.645 ;
        RECT  10.735 1.935 11.230 2.235 ;
        RECT  10.965 2.480 11.195 3.300 ;
        RECT  10.985 1.280 11.040 1.620 ;
        RECT  10.505 1.310 10.735 3.845 ;
        RECT  9.765 1.310 10.505 1.540 ;
        RECT  9.530 2.975 10.505 3.205 ;
        RECT  9.920 2.255 10.235 2.485 ;
        RECT  9.690 1.775 9.920 2.485 ;
        RECT  9.605 1.200 9.765 1.540 ;
        RECT  8.460 1.775 9.690 2.005 ;
        RECT  9.425 0.630 9.605 1.540 ;
        RECT  9.375 0.630 9.425 1.485 ;
        RECT  9.070 2.240 9.410 2.580 ;
        RECT  9.265 0.630 9.375 0.970 ;
        RECT  8.885 2.350 9.070 2.580 ;
        RECT  8.655 2.350 8.885 3.845 ;
        RECT  6.295 3.615 8.655 3.845 ;
        RECT  8.425 1.300 8.460 2.005 ;
        RECT  8.195 1.300 8.425 3.325 ;
        RECT  8.120 1.300 8.195 1.640 ;
        RECT  6.820 3.095 8.195 3.325 ;
        RECT  7.735 2.005 7.965 2.380 ;
        RECT  6.080 2.005 7.735 2.235 ;
        RECT  6.590 2.525 6.820 3.325 ;
        RECT  6.385 2.525 6.590 2.755 ;
        RECT  6.065 3.615 6.295 4.345 ;
        RECT  5.885 1.010 6.080 2.735 ;
        RECT  5.340 4.115 6.065 4.345 ;
        RECT  5.850 0.955 5.885 2.735 ;
        RECT  5.545 0.955 5.850 1.295 ;
        RECT  5.800 2.505 5.850 2.735 ;
        RECT  5.570 2.505 5.800 3.800 ;
        RECT  5.340 1.770 5.605 2.110 ;
        RECT  5.265 1.770 5.340 4.345 ;
        RECT  5.110 1.825 5.265 4.345 ;
        RECT  3.500 4.115 5.110 4.345 ;
        RECT  3.935 0.710 5.085 0.940 ;
        RECT  3.960 3.570 4.865 3.800 ;
        RECT  4.415 2.580 4.420 3.150 ;
        RECT  4.190 1.355 4.415 3.150 ;
        RECT  4.185 1.355 4.190 2.810 ;
        RECT  2.735 1.870 4.185 2.100 ;
        RECT  3.730 3.055 3.960 3.800 ;
        RECT  3.705 0.710 3.935 1.640 ;
        RECT  2.100 3.055 3.730 3.285 ;
        RECT  2.100 1.410 3.705 1.640 ;
        RECT  3.270 3.515 3.500 4.345 ;
        RECT  0.520 3.515 3.270 3.745 ;
        RECT  2.395 1.870 2.735 2.690 ;
        RECT  1.860 1.870 2.395 2.100 ;
        RECT  1.630 0.685 1.860 2.100 ;
        RECT  1.390 0.685 1.630 0.915 ;
        RECT  0.410 1.420 0.520 1.760 ;
        RECT  0.410 2.870 0.520 3.745 ;
        RECT  0.290 1.420 0.410 3.745 ;
        RECT  0.180 1.420 0.290 3.210 ;
    END
END SDFFSRHQX1

MACRO SDFFSRXL
    CLASS CORE ;
    FOREIGN SDFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 4.035 14.010 4.265 ;
        RECT  13.415 4.035 13.645 4.365 ;
        RECT  11.000 4.135 13.415 4.365 ;
        RECT  10.770 4.125 11.000 4.365 ;
        RECT  8.375 4.125 10.770 4.355 ;
        RECT  8.145 4.005 8.375 4.355 ;
        RECT  7.320 4.005 8.145 4.235 ;
        RECT  7.090 4.005 7.320 4.365 ;
        RECT  7.045 4.085 7.090 4.365 ;
        RECT  6.820 4.135 7.045 4.365 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.230 2.165 3.505 2.505 ;
        RECT  3.165 2.165 3.230 3.195 ;
        RECT  3.000 2.220 3.165 3.195 ;
        RECT  2.855 2.965 3.000 3.195 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.235 0.670 1.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.800 1.785 9.025 2.175 ;
        RECT  8.675 1.765 8.800 2.175 ;
        RECT  8.485 1.765 8.675 2.155 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 1.340 17.640 1.845 ;
        RECT  17.430 1.285 17.605 1.845 ;
        RECT  17.280 1.285 17.430 3.400 ;
        RECT  17.200 1.285 17.280 3.455 ;
        RECT  16.940 3.115 17.200 3.455 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.925 1.340 18.960 1.845 ;
        RECT  18.695 1.340 18.925 3.525 ;
        RECT  18.620 1.340 18.695 1.845 ;
        RECT  18.300 3.220 18.695 3.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.380 2.500 2.730 ;
        RECT  2.240 2.335 2.425 2.730 ;
        RECT  1.900 2.280 2.240 2.730 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  10.290 2.250 11.080 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.490 -0.400 19.140 0.400 ;
        RECT  18.150 -0.400 18.490 0.575 ;
        RECT  16.930 -0.400 18.150 0.400 ;
        RECT  16.590 -0.400 16.930 0.575 ;
        RECT  13.735 -0.400 16.590 0.400 ;
        RECT  13.395 -0.400 13.735 0.575 ;
        RECT  11.170 -0.400 13.395 0.400 ;
        RECT  10.830 -0.400 11.170 1.485 ;
        RECT  9.395 -0.400 10.830 0.400 ;
        RECT  9.165 -0.400 9.395 0.900 ;
        RECT  6.475 -0.400 9.165 0.400 ;
        RECT  6.135 -0.400 6.475 0.900 ;
        RECT  3.710 -0.400 6.135 0.400 ;
        RECT  3.370 -0.400 3.710 0.575 ;
        RECT  1.380 -0.400 3.370 0.400 ;
        RECT  1.040 -0.400 1.380 0.920 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.880 4.640 19.140 5.440 ;
        RECT  17.540 4.465 17.880 5.440 ;
        RECT  15.850 4.640 17.540 5.440 ;
        RECT  15.510 3.395 15.850 5.440 ;
        RECT  14.685 4.640 15.510 5.440 ;
        RECT  14.455 3.395 14.685 5.440 ;
        RECT  13.770 3.395 14.455 3.625 ;
        RECT  7.915 4.640 14.455 5.440 ;
        RECT  13.410 3.310 13.770 3.625 ;
        RECT  13.185 3.395 13.410 3.625 ;
        RECT  12.955 3.395 13.185 3.845 ;
        RECT  11.500 3.615 12.955 3.845 ;
        RECT  11.270 3.570 11.500 3.845 ;
        RECT  11.075 3.570 11.270 3.800 ;
        RECT  10.735 3.460 11.075 3.800 ;
        RECT  7.575 4.465 7.915 5.440 ;
        RECT  6.590 4.640 7.575 5.440 ;
        RECT  6.250 4.465 6.590 5.440 ;
        RECT  3.480 4.640 6.250 5.440 ;
        RECT  3.140 4.465 3.480 5.440 ;
        RECT  0.890 4.640 3.140 5.440 ;
        RECT  0.550 4.465 0.890 5.440 ;
        RECT  0.000 4.640 0.550 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.935 2.330 18.275 2.670 ;
        RECT  17.905 2.440 17.935 2.670 ;
        RECT  17.675 2.440 17.905 3.995 ;
        RECT  16.595 3.765 17.675 3.995 ;
        RECT  16.600 1.170 16.940 1.510 ;
        RECT  16.595 1.280 16.600 1.510 ;
        RECT  16.365 1.280 16.595 3.995 ;
        RECT  16.230 3.395 16.365 3.735 ;
        RECT  15.885 0.980 16.135 1.320 ;
        RECT  16.080 2.065 16.135 2.405 ;
        RECT  16.025 2.065 16.080 3.165 ;
        RECT  15.850 1.825 16.025 3.165 ;
        RECT  15.655 0.630 15.885 1.320 ;
        RECT  15.795 1.825 15.850 2.405 ;
        RECT  14.290 2.935 15.850 3.165 ;
        RECT  15.425 1.825 15.795 2.055 ;
        RECT  14.535 0.630 15.655 0.860 ;
        RECT  15.195 1.090 15.425 2.055 ;
        RECT  14.995 1.090 15.195 1.320 ;
        RECT  14.470 1.855 14.700 2.230 ;
        RECT  14.305 0.630 14.535 1.290 ;
        RECT  13.345 1.855 14.470 2.085 ;
        RECT  14.195 0.950 14.305 1.290 ;
        RECT  14.060 2.670 14.290 3.165 ;
        RECT  13.575 2.670 14.060 2.900 ;
        RECT  13.235 2.560 13.575 2.900 ;
        RECT  13.115 1.250 13.345 2.085 ;
        RECT  12.695 1.250 13.115 1.480 ;
        RECT  11.825 0.720 12.985 0.950 ;
        RECT  12.465 1.250 12.695 3.360 ;
        RECT  12.395 1.250 12.465 1.535 ;
        RECT  12.055 3.130 12.465 3.360 ;
        RECT  12.165 1.195 12.395 1.535 ;
        RECT  11.825 2.430 12.150 2.770 ;
        RECT  11.595 0.720 11.825 3.125 ;
        RECT  10.315 1.745 11.595 1.975 ;
        RECT  10.300 2.895 11.595 3.125 ;
        RECT  10.085 1.370 10.315 1.975 ;
        RECT  10.070 2.895 10.300 3.835 ;
        RECT  9.855 0.740 10.215 0.970 ;
        RECT  8.835 3.605 10.070 3.835 ;
        RECT  9.625 0.740 9.855 1.365 ;
        RECT  7.950 1.135 9.625 1.365 ;
        RECT  9.525 1.635 9.580 3.030 ;
        RECT  9.350 1.635 9.525 3.375 ;
        RECT  9.200 2.460 9.350 3.375 ;
        RECT  9.150 2.800 9.200 3.375 ;
        RECT  9.065 2.905 9.150 3.375 ;
        RECT  8.380 2.905 9.065 3.135 ;
        RECT  8.605 3.545 8.835 3.835 ;
        RECT  6.000 3.545 8.605 3.775 ;
        RECT  8.150 2.540 8.380 3.135 ;
        RECT  7.920 1.120 7.950 1.460 ;
        RECT  7.690 1.120 7.920 3.135 ;
        RECT  7.610 1.120 7.690 1.460 ;
        RECT  7.370 2.905 7.690 3.135 ;
        RECT  7.215 1.840 7.445 2.205 ;
        RECT  6.325 2.905 7.370 3.260 ;
        RECT  5.865 1.975 7.215 2.205 ;
        RECT  6.095 2.510 6.325 3.260 ;
        RECT  5.770 3.545 6.000 4.365 ;
        RECT  5.635 0.955 5.865 2.965 ;
        RECT  5.420 4.135 5.770 4.365 ;
        RECT  5.310 0.955 5.635 1.240 ;
        RECT  5.335 2.735 5.635 2.965 ;
        RECT  5.175 1.770 5.405 2.225 ;
        RECT  5.105 2.735 5.335 3.820 ;
        RECT  4.970 0.900 5.310 1.240 ;
        RECT  4.710 1.995 5.175 2.225 ;
        RECT  4.710 3.280 4.785 3.645 ;
        RECT  4.510 1.485 4.710 3.645 ;
        RECT  4.480 1.430 4.510 3.645 ;
        RECT  4.330 0.745 4.505 0.975 ;
        RECT  4.170 1.430 4.480 1.770 ;
        RECT  3.835 3.145 4.480 3.485 ;
        RECT  4.100 0.745 4.330 1.095 ;
        RECT  4.075 3.945 4.305 4.320 ;
        RECT  2.860 0.865 4.100 1.095 ;
        RECT  3.255 3.945 4.075 4.175 ;
        RECT  3.025 3.615 3.255 4.175 ;
        RECT  2.295 3.615 3.025 3.845 ;
        RECT  2.630 0.865 2.860 1.585 ;
        RECT  2.490 1.355 2.630 1.585 ;
        RECT  1.775 4.145 2.535 4.375 ;
        RECT  2.260 1.355 2.490 1.960 ;
        RECT  2.065 3.300 2.295 3.845 ;
        RECT  2.005 0.675 2.185 0.905 ;
        RECT  1.955 3.300 2.065 3.640 ;
        RECT  1.775 0.675 2.005 1.625 ;
        RECT  1.570 1.395 1.775 1.625 ;
        RECT  1.455 4.145 1.775 4.410 ;
        RECT  1.340 1.395 1.570 2.590 ;
        RECT  1.225 3.945 1.455 4.410 ;
        RECT  1.335 2.255 1.340 2.590 ;
        RECT  0.995 2.255 1.335 2.645 ;
        RECT  0.455 3.945 1.225 4.175 ;
        RECT  0.455 2.255 0.995 2.485 ;
        RECT  0.225 2.255 0.455 4.175 ;
    END
END SDFFSRXL

MACRO SDFFSRX4
    CLASS CORE ;
    FOREIGN SDFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRXL ;
    SIZE 25.740 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 4.000 16.960 4.230 ;
        RECT  11.140 4.000 11.370 4.290 ;
        RECT  11.005 4.060 11.140 4.290 ;
        RECT  10.775 4.060 11.005 4.335 ;
        RECT  7.300 4.105 10.775 4.335 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 2.180 3.085 3.195 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 2.405 1.205 2.835 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.235 2.295 9.705 2.790 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.620 1.420 23.640 1.845 ;
        RECT  23.620 2.635 23.640 3.195 ;
        RECT  23.300 1.420 23.620 3.220 ;
        RECT  23.240 1.820 23.300 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.920 1.820 24.940 3.220 ;
        RECT  24.580 1.420 24.920 3.220 ;
        RECT  24.560 1.820 24.580 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 2.405 2.425 2.815 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.880 4.060 2.265 ;
        RECT  3.515 1.845 3.745 2.265 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.560 -0.400 25.740 0.400 ;
        RECT  25.220 -0.400 25.560 1.030 ;
        RECT  24.280 -0.400 25.220 0.400 ;
        RECT  23.940 -0.400 24.280 1.045 ;
        RECT  22.960 -0.400 23.940 0.400 ;
        RECT  22.620 -0.400 22.960 0.575 ;
        RECT  17.790 -0.400 22.620 0.400 ;
        RECT  17.450 -0.400 17.790 1.050 ;
        RECT  14.850 -0.400 17.450 0.400 ;
        RECT  14.620 -0.400 14.850 1.145 ;
        RECT  12.305 -0.400 14.620 0.400 ;
        RECT  11.965 -0.400 12.305 1.640 ;
        RECT  9.645 -0.400 11.965 0.400 ;
        RECT  9.415 -0.400 9.645 0.875 ;
        RECT  6.975 -0.400 9.415 0.400 ;
        RECT  6.635 -0.400 6.975 0.845 ;
        RECT  3.670 -0.400 6.635 0.400 ;
        RECT  3.330 -0.400 3.670 0.575 ;
        RECT  1.170 -0.400 3.330 0.400 ;
        RECT  0.830 -0.400 1.170 0.900 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.560 4.640 25.740 5.440 ;
        RECT  25.220 4.035 25.560 5.440 ;
        RECT  24.280 4.640 25.220 5.440 ;
        RECT  23.940 4.035 24.280 5.440 ;
        RECT  23.000 4.640 23.940 5.440 ;
        RECT  22.660 4.035 23.000 5.440 ;
        RECT  20.250 4.640 22.660 5.440 ;
        RECT  19.910 3.300 20.250 5.440 ;
        RECT  18.190 4.640 19.910 5.440 ;
        RECT  17.960 2.920 18.190 5.440 ;
        RECT  15.985 4.640 17.960 5.440 ;
        RECT  15.645 4.465 15.985 5.440 ;
        RECT  14.830 4.640 15.645 5.440 ;
        RECT  14.490 4.465 14.830 5.440 ;
        RECT  12.165 4.640 14.490 5.440 ;
        RECT  11.825 4.465 12.165 5.440 ;
        RECT  7.050 4.640 11.825 5.440 ;
        RECT  6.710 4.465 7.050 5.440 ;
        RECT  3.525 4.640 6.710 5.440 ;
        RECT  3.185 4.465 3.525 5.440 ;
        RECT  1.140 4.640 3.185 5.440 ;
        RECT  0.800 4.465 1.140 5.440 ;
        RECT  0.000 4.640 0.800 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  25.455 2.210 25.510 2.550 ;
        RECT  25.225 2.210 25.455 3.740 ;
        RECT  25.170 2.210 25.225 2.550 ;
        RECT  22.935 3.510 25.225 3.740 ;
        RECT  22.705 1.670 22.935 3.740 ;
        RECT  22.040 1.670 22.705 1.900 ;
        RECT  22.240 3.400 22.705 3.740 ;
        RECT  21.575 2.160 22.390 2.500 ;
        RECT  21.900 3.165 22.240 3.975 ;
        RECT  21.810 1.440 22.040 1.900 ;
        RECT  21.540 1.375 21.575 3.015 ;
        RECT  21.345 1.375 21.540 3.845 ;
        RECT  21.125 0.675 21.355 1.030 ;
        RECT  20.690 1.375 21.345 1.605 ;
        RECT  21.310 2.785 21.345 3.845 ;
        RECT  21.200 2.840 21.310 3.845 ;
        RECT  18.970 2.840 21.200 3.070 ;
        RECT  19.970 0.675 21.125 0.905 ;
        RECT  20.885 1.860 21.115 2.260 ;
        RECT  18.750 1.860 20.885 2.090 ;
        RECT  20.320 1.205 20.690 1.605 ;
        RECT  19.345 1.375 20.320 1.605 ;
        RECT  19.630 0.675 19.970 1.050 ;
        RECT  18.515 0.675 19.630 0.905 ;
        RECT  19.115 1.140 19.345 1.605 ;
        RECT  18.905 1.140 19.115 1.370 ;
        RECT  18.860 2.840 18.970 3.835 ;
        RECT  18.630 2.455 18.860 3.835 ;
        RECT  18.465 1.860 18.750 2.155 ;
        RECT  17.470 2.455 18.630 2.685 ;
        RECT  18.405 0.675 18.515 1.290 ;
        RECT  16.320 1.925 18.465 2.155 ;
        RECT  18.285 0.675 18.405 1.605 ;
        RECT  18.175 0.950 18.285 1.605 ;
        RECT  17.015 1.375 18.175 1.605 ;
        RECT  17.395 3.535 17.625 4.410 ;
        RECT  17.240 2.455 17.470 3.305 ;
        RECT  10.835 3.535 17.395 3.765 ;
        RECT  15.395 3.075 17.240 3.305 ;
        RECT  16.785 0.970 17.015 1.605 ;
        RECT  16.090 0.865 16.320 2.155 ;
        RECT  15.925 0.865 16.090 1.095 ;
        RECT  15.930 1.925 16.090 2.155 ;
        RECT  15.930 2.505 15.985 2.845 ;
        RECT  15.700 1.925 15.930 2.845 ;
        RECT  14.160 1.405 15.860 1.635 ;
        RECT  13.695 1.925 15.700 2.155 ;
        RECT  15.645 2.505 15.700 2.845 ;
        RECT  15.165 2.385 15.395 3.305 ;
        RECT  14.960 2.385 15.165 2.615 ;
        RECT  13.930 0.675 14.160 1.635 ;
        RECT  12.895 0.675 13.930 0.905 ;
        RECT  13.530 1.755 13.695 3.135 ;
        RECT  13.495 1.220 13.530 3.135 ;
        RECT  13.465 1.220 13.495 3.190 ;
        RECT  13.300 1.220 13.465 1.985 ;
        RECT  13.155 2.850 13.465 3.190 ;
        RECT  12.895 2.275 13.230 2.505 ;
        RECT  12.665 0.675 12.895 2.505 ;
        RECT  11.335 2.045 12.665 2.275 ;
        RECT  11.205 1.400 11.545 1.740 ;
        RECT  11.300 2.910 11.545 3.250 ;
        RECT  10.110 0.740 11.355 0.970 ;
        RECT  11.205 2.565 11.300 3.250 ;
        RECT  11.040 1.455 11.205 1.740 ;
        RECT  11.070 2.565 11.205 3.195 ;
        RECT  11.040 2.565 11.070 2.795 ;
        RECT  10.810 1.455 11.040 2.795 ;
        RECT  10.605 3.085 10.835 3.765 ;
        RECT  10.585 2.165 10.810 2.505 ;
        RECT  10.245 3.085 10.605 3.315 ;
        RECT  10.245 1.570 10.395 1.910 ;
        RECT  10.320 3.605 10.375 3.835 ;
        RECT  10.090 3.605 10.320 3.840 ;
        RECT  10.055 1.570 10.245 3.315 ;
        RECT  9.880 0.740 10.110 1.335 ;
        RECT  6.325 3.610 10.090 3.840 ;
        RECT  10.015 1.625 10.055 3.315 ;
        RECT  8.810 3.085 10.015 3.315 ;
        RECT  8.340 1.105 9.880 1.335 ;
        RECT  8.580 2.280 8.810 3.315 ;
        RECT  8.110 1.105 8.340 3.375 ;
        RECT  8.040 1.105 8.110 1.435 ;
        RECT  6.705 3.145 8.110 3.375 ;
        RECT  7.645 1.775 7.875 2.240 ;
        RECT  5.865 1.775 7.645 2.005 ;
        RECT  6.705 2.330 6.760 2.670 ;
        RECT  6.475 2.330 6.705 3.375 ;
        RECT  6.420 2.330 6.475 2.670 ;
        RECT  6.095 3.610 6.325 4.410 ;
        RECT  5.230 4.180 6.095 4.410 ;
        RECT  5.795 0.665 5.865 2.005 ;
        RECT  5.690 0.665 5.795 2.415 ;
        RECT  5.565 0.665 5.690 3.805 ;
        RECT  5.420 0.665 5.565 0.895 ;
        RECT  5.460 2.185 5.565 3.805 ;
        RECT  4.615 1.520 5.250 1.860 ;
        RECT  5.000 3.130 5.230 4.410 ;
        RECT  4.805 0.675 5.035 0.905 ;
        RECT  4.615 3.130 5.000 3.360 ;
        RECT  4.575 0.675 4.805 1.095 ;
        RECT  4.540 3.735 4.770 4.100 ;
        RECT  4.385 1.415 4.615 3.360 ;
        RECT  2.605 0.865 4.575 1.095 ;
        RECT  3.585 3.735 4.540 3.965 ;
        RECT  4.205 1.415 4.385 1.645 ;
        RECT  3.945 3.020 4.385 3.360 ;
        RECT  3.355 3.605 3.585 3.965 ;
        RECT  2.400 3.605 3.355 3.835 ;
        RECT  1.685 4.125 2.750 4.355 ;
        RECT  2.500 0.865 2.605 1.545 ;
        RECT  2.375 0.865 2.500 1.600 ;
        RECT  2.170 3.130 2.400 3.835 ;
        RECT  2.160 1.260 2.375 1.600 ;
        RECT  2.060 3.130 2.170 3.470 ;
        RECT  1.455 3.185 1.685 4.355 ;
        RECT  0.520 1.865 1.560 2.095 ;
        RECT  0.520 3.185 1.455 3.415 ;
        RECT  0.405 1.400 0.520 2.095 ;
        RECT  0.405 3.130 0.520 3.470 ;
        RECT  0.180 1.400 0.405 3.470 ;
        RECT  0.175 1.400 0.180 3.415 ;
    END
END SDFFSRX4

MACRO SDFFSRX2
    CLASS CORE ;
    FOREIGN SDFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 4.035 14.010 4.265 ;
        RECT  13.415 4.035 13.645 4.365 ;
        RECT  11.000 4.135 13.415 4.365 ;
        RECT  10.770 4.125 11.000 4.365 ;
        RECT  8.375 4.125 10.770 4.355 ;
        RECT  8.145 4.005 8.375 4.355 ;
        RECT  7.320 4.005 8.145 4.235 ;
        RECT  7.090 4.005 7.320 4.365 ;
        RECT  7.045 4.085 7.090 4.365 ;
        RECT  6.820 4.135 7.045 4.365 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.230 2.200 3.340 2.540 ;
        RECT  3.000 2.200 3.230 3.195 ;
        RECT  2.855 2.965 3.000 3.195 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.690 2.820 1.180 3.340 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.465 1.785 9.025 2.175 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.595 1.845 17.605 2.075 ;
        RECT  17.300 1.325 17.595 2.100 ;
        RECT  17.300 2.915 17.355 3.255 ;
        RECT  17.255 1.325 17.300 3.255 ;
        RECT  17.070 1.845 17.255 3.255 ;
        RECT  17.015 2.915 17.070 3.255 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.925 2.940 19.000 3.220 ;
        RECT  18.875 1.380 18.925 3.220 ;
        RECT  18.695 1.325 18.875 3.220 ;
        RECT  18.535 1.325 18.695 1.665 ;
        RECT  18.295 2.915 18.695 3.255 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.380 2.500 2.730 ;
        RECT  2.240 2.335 2.425 2.730 ;
        RECT  1.900 2.280 2.240 2.730 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  10.290 2.250 11.080 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.235 -0.400 19.140 0.400 ;
        RECT  17.895 -0.400 18.235 0.950 ;
        RECT  16.815 -0.400 17.895 0.400 ;
        RECT  16.455 -0.400 16.815 0.575 ;
        RECT  13.755 -0.400 16.455 0.400 ;
        RECT  13.415 -0.400 13.755 0.575 ;
        RECT  11.170 -0.400 13.415 0.400 ;
        RECT  10.830 -0.400 11.170 1.400 ;
        RECT  9.435 -0.400 10.830 0.400 ;
        RECT  9.205 -0.400 9.435 0.900 ;
        RECT  6.475 -0.400 9.205 0.400 ;
        RECT  6.135 -0.400 6.475 0.900 ;
        RECT  3.710 -0.400 6.135 0.400 ;
        RECT  3.370 -0.400 3.710 0.575 ;
        RECT  1.380 -0.400 3.370 0.400 ;
        RECT  1.040 -0.400 1.380 0.920 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.995 4.640 19.140 5.440 ;
        RECT  17.655 4.065 17.995 5.440 ;
        RECT  15.770 4.640 17.655 5.440 ;
        RECT  15.430 3.560 15.770 5.440 ;
        RECT  14.685 4.640 15.430 5.440 ;
        RECT  14.455 3.485 14.685 5.440 ;
        RECT  13.185 3.485 14.455 3.715 ;
        RECT  7.915 4.640 14.455 5.440 ;
        RECT  12.955 3.485 13.185 3.845 ;
        RECT  11.245 3.615 12.955 3.845 ;
        RECT  11.015 3.515 11.245 3.845 ;
        RECT  10.775 3.515 11.015 3.745 ;
        RECT  7.575 4.465 7.915 5.440 ;
        RECT  6.590 4.640 7.575 5.440 ;
        RECT  6.250 4.465 6.590 5.440 ;
        RECT  3.480 4.640 6.250 5.440 ;
        RECT  3.140 4.465 3.480 5.440 ;
        RECT  0.890 4.640 3.140 5.440 ;
        RECT  0.550 4.465 0.890 5.440 ;
        RECT  0.000 4.640 0.550 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.235 2.085 18.465 2.675 ;
        RECT  17.960 2.445 18.235 2.675 ;
        RECT  17.730 2.445 17.960 3.830 ;
        RECT  16.555 3.600 17.730 3.830 ;
        RECT  16.555 1.170 16.815 1.510 ;
        RECT  16.475 1.170 16.555 4.005 ;
        RECT  16.325 1.225 16.475 4.005 ;
        RECT  16.155 3.665 16.325 4.005 ;
        RECT  15.860 1.825 16.090 3.165 ;
        RECT  15.655 0.700 15.995 1.510 ;
        RECT  15.300 1.825 15.860 2.055 ;
        RECT  14.095 2.935 15.860 3.165 ;
        RECT  14.555 0.745 15.655 0.975 ;
        RECT  15.070 1.275 15.300 2.055 ;
        RECT  14.935 1.275 15.070 1.505 ;
        RECT  14.470 1.855 14.700 2.230 ;
        RECT  14.215 0.740 14.555 1.550 ;
        RECT  13.345 1.855 14.470 2.085 ;
        RECT  13.865 2.615 14.095 3.165 ;
        RECT  13.010 2.615 13.865 2.845 ;
        RECT  13.115 1.335 13.345 2.085 ;
        RECT  12.695 1.335 13.115 1.565 ;
        RECT  11.820 0.735 12.985 0.965 ;
        RECT  12.465 1.335 12.695 3.325 ;
        RECT  12.450 1.335 12.465 1.620 ;
        RECT  12.055 3.095 12.465 3.325 ;
        RECT  12.110 1.280 12.450 1.620 ;
        RECT  11.840 2.525 12.150 2.755 ;
        RECT  11.820 1.745 11.840 2.755 ;
        RECT  11.590 0.735 11.820 3.225 ;
        RECT  10.355 1.745 11.590 1.975 ;
        RECT  10.340 2.995 11.590 3.225 ;
        RECT  10.125 1.370 10.355 1.975 ;
        RECT  10.110 2.995 10.340 3.835 ;
        RECT  9.895 0.735 10.215 0.965 ;
        RECT  8.835 3.605 10.110 3.835 ;
        RECT  9.665 0.735 9.895 1.365 ;
        RECT  9.585 2.460 9.675 2.800 ;
        RECT  7.950 1.135 9.665 1.365 ;
        RECT  9.355 1.600 9.585 3.375 ;
        RECT  9.335 2.460 9.355 3.375 ;
        RECT  9.295 2.515 9.335 3.375 ;
        RECT  9.065 2.905 9.295 3.375 ;
        RECT  8.380 2.905 9.065 3.135 ;
        RECT  8.605 3.545 8.835 3.835 ;
        RECT  6.000 3.545 8.605 3.775 ;
        RECT  8.150 2.540 8.380 3.135 ;
        RECT  7.920 1.120 7.950 1.460 ;
        RECT  7.690 1.120 7.920 3.135 ;
        RECT  7.610 1.120 7.690 1.460 ;
        RECT  7.370 2.905 7.690 3.135 ;
        RECT  7.215 1.840 7.445 2.205 ;
        RECT  6.325 2.905 7.370 3.260 ;
        RECT  5.865 1.975 7.215 2.205 ;
        RECT  6.095 2.510 6.325 3.260 ;
        RECT  5.770 3.545 6.000 4.365 ;
        RECT  5.635 0.955 5.865 2.965 ;
        RECT  5.420 4.135 5.770 4.365 ;
        RECT  5.310 0.955 5.635 1.240 ;
        RECT  5.335 2.735 5.635 2.965 ;
        RECT  5.175 1.770 5.405 2.225 ;
        RECT  5.105 2.735 5.335 3.820 ;
        RECT  4.970 0.900 5.310 1.240 ;
        RECT  4.710 1.995 5.175 2.225 ;
        RECT  4.710 3.280 4.785 3.645 ;
        RECT  4.510 1.455 4.710 3.645 ;
        RECT  4.495 1.400 4.510 3.645 ;
        RECT  4.290 0.695 4.505 0.925 ;
        RECT  4.480 1.400 4.495 3.535 ;
        RECT  4.170 1.400 4.480 1.740 ;
        RECT  3.835 3.250 4.480 3.535 ;
        RECT  4.075 3.945 4.305 4.320 ;
        RECT  4.060 0.695 4.290 1.095 ;
        RECT  3.255 3.945 4.075 4.175 ;
        RECT  2.860 0.865 4.060 1.095 ;
        RECT  3.025 3.615 3.255 4.175 ;
        RECT  2.295 3.615 3.025 3.845 ;
        RECT  2.630 0.865 2.860 1.585 ;
        RECT  2.490 1.355 2.630 1.585 ;
        RECT  1.455 4.145 2.535 4.375 ;
        RECT  2.260 1.355 2.490 1.960 ;
        RECT  2.065 3.300 2.295 3.845 ;
        RECT  2.005 0.675 2.185 0.905 ;
        RECT  1.955 3.300 2.065 3.640 ;
        RECT  1.775 0.675 2.005 1.625 ;
        RECT  1.570 1.395 1.775 1.625 ;
        RECT  1.340 1.395 1.570 2.490 ;
        RECT  1.225 3.945 1.455 4.375 ;
        RECT  1.230 2.150 1.340 2.490 ;
        RECT  0.455 2.255 1.230 2.485 ;
        RECT  0.455 3.945 1.225 4.175 ;
        RECT  0.225 2.255 0.455 4.175 ;
    END
END SDFFSRX2

MACRO SDFFSRX1
    CLASS CORE ;
    FOREIGN SDFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 4.035 14.010 4.265 ;
        RECT  13.415 4.035 13.645 4.365 ;
        RECT  11.000 4.135 13.415 4.365 ;
        RECT  10.770 4.125 11.000 4.365 ;
        RECT  8.375 4.125 10.770 4.355 ;
        RECT  8.145 4.005 8.375 4.355 ;
        RECT  7.320 4.005 8.145 4.235 ;
        RECT  7.090 4.005 7.320 4.365 ;
        RECT  7.045 4.085 7.090 4.365 ;
        RECT  6.820 4.135 7.045 4.365 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.230 2.200 3.340 2.540 ;
        RECT  3.000 2.200 3.230 3.195 ;
        RECT  2.855 2.965 3.000 3.195 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.690 2.820 1.180 3.340 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.485 1.785 9.025 2.175 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.615 1.095 17.770 1.435 ;
        RECT  17.605 1.095 17.615 3.205 ;
        RECT  17.385 1.095 17.605 3.400 ;
        RECT  17.155 2.965 17.385 3.400 ;
        RECT  17.100 3.170 17.155 3.400 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.170 1.050 19.315 3.185 ;
        RECT  19.085 1.050 19.170 3.780 ;
        RECT  18.950 1.050 19.085 1.390 ;
        RECT  19.000 2.940 19.085 3.780 ;
        RECT  18.830 2.955 19.000 3.780 ;
        RECT  18.695 2.955 18.830 3.195 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.380 2.500 2.730 ;
        RECT  2.240 2.335 2.425 2.730 ;
        RECT  1.900 2.280 2.240 2.730 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  10.290 2.250 11.080 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.530 -0.400 19.800 0.400 ;
        RECT  18.190 -0.400 18.530 1.390 ;
        RECT  16.795 -0.400 18.190 0.400 ;
        RECT  16.455 -0.400 16.795 0.575 ;
        RECT  13.755 -0.400 16.455 0.400 ;
        RECT  13.415 -0.400 13.755 0.575 ;
        RECT  11.170 -0.400 13.415 0.400 ;
        RECT  10.830 -0.400 11.170 1.485 ;
        RECT  9.395 -0.400 10.830 0.400 ;
        RECT  9.165 -0.400 9.395 0.900 ;
        RECT  6.475 -0.400 9.165 0.400 ;
        RECT  6.135 -0.400 6.475 0.900 ;
        RECT  3.710 -0.400 6.135 0.400 ;
        RECT  3.370 -0.400 3.710 0.575 ;
        RECT  1.380 -0.400 3.370 0.400 ;
        RECT  1.040 -0.400 1.380 0.920 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.350 4.640 19.800 5.440 ;
        RECT  18.010 4.090 18.350 5.440 ;
        RECT  15.850 4.640 18.010 5.440 ;
        RECT  15.510 3.395 15.850 5.440 ;
        RECT  14.685 4.640 15.510 5.440 ;
        RECT  14.455 3.430 14.685 5.440 ;
        RECT  13.185 3.430 14.455 3.660 ;
        RECT  7.915 4.640 14.455 5.440 ;
        RECT  12.955 3.430 13.185 3.845 ;
        RECT  11.245 3.615 12.955 3.845 ;
        RECT  11.075 3.455 11.245 3.845 ;
        RECT  11.015 3.400 11.075 3.845 ;
        RECT  10.735 3.400 11.015 3.740 ;
        RECT  7.575 4.465 7.915 5.440 ;
        RECT  6.590 4.640 7.575 5.440 ;
        RECT  6.250 4.465 6.590 5.440 ;
        RECT  3.480 4.640 6.250 5.440 ;
        RECT  3.140 4.465 3.480 5.440 ;
        RECT  0.890 4.640 3.140 5.440 ;
        RECT  0.550 4.465 0.890 5.440 ;
        RECT  0.000 4.640 0.550 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.260 2.145 18.730 2.375 ;
        RECT  18.030 2.145 18.260 3.860 ;
        RECT  16.865 3.630 18.030 3.860 ;
        RECT  16.815 1.225 16.865 3.860 ;
        RECT  16.635 1.170 16.815 3.860 ;
        RECT  16.475 1.170 16.635 1.510 ;
        RECT  16.230 3.395 16.635 3.735 ;
        RECT  16.220 2.300 16.330 2.640 ;
        RECT  15.990 1.825 16.220 3.165 ;
        RECT  15.885 0.980 15.995 1.320 ;
        RECT  15.300 1.825 15.990 2.055 ;
        RECT  14.095 2.935 15.990 3.165 ;
        RECT  15.655 0.630 15.885 1.320 ;
        RECT  14.555 0.630 15.655 0.860 ;
        RECT  15.070 1.090 15.300 2.055 ;
        RECT  14.935 1.090 15.070 1.320 ;
        RECT  14.470 1.855 14.700 2.230 ;
        RECT  14.325 0.630 14.555 1.290 ;
        RECT  13.345 1.855 14.470 2.085 ;
        RECT  14.215 0.950 14.325 1.290 ;
        RECT  13.865 2.615 14.095 3.165 ;
        RECT  13.010 2.615 13.865 2.845 ;
        RECT  13.115 1.250 13.345 2.085 ;
        RECT  12.695 1.250 13.115 1.480 ;
        RECT  11.820 0.735 12.985 0.965 ;
        RECT  12.465 1.250 12.695 3.330 ;
        RECT  12.450 1.250 12.465 1.535 ;
        RECT  12.055 3.100 12.465 3.330 ;
        RECT  12.110 1.195 12.450 1.535 ;
        RECT  11.840 2.525 12.150 2.755 ;
        RECT  11.820 1.745 11.840 2.755 ;
        RECT  11.590 0.735 11.820 3.125 ;
        RECT  10.315 1.745 11.590 1.975 ;
        RECT  10.300 2.895 11.590 3.125 ;
        RECT  10.085 1.370 10.315 1.975 ;
        RECT  10.070 2.895 10.300 3.835 ;
        RECT  9.855 0.740 10.215 0.970 ;
        RECT  8.835 3.605 10.070 3.835 ;
        RECT  9.625 0.740 9.855 1.365 ;
        RECT  9.580 2.460 9.675 2.800 ;
        RECT  7.950 1.135 9.625 1.365 ;
        RECT  9.350 1.635 9.580 3.375 ;
        RECT  9.335 2.460 9.350 3.375 ;
        RECT  9.295 2.515 9.335 3.375 ;
        RECT  9.065 2.905 9.295 3.375 ;
        RECT  8.380 2.905 9.065 3.135 ;
        RECT  8.605 3.545 8.835 3.835 ;
        RECT  6.000 3.545 8.605 3.775 ;
        RECT  8.150 2.540 8.380 3.135 ;
        RECT  7.920 1.120 7.950 1.460 ;
        RECT  7.690 1.120 7.920 3.135 ;
        RECT  7.610 1.120 7.690 1.460 ;
        RECT  7.370 2.905 7.690 3.135 ;
        RECT  7.215 1.840 7.445 2.205 ;
        RECT  6.325 2.905 7.370 3.260 ;
        RECT  5.865 1.975 7.215 2.205 ;
        RECT  6.095 2.510 6.325 3.260 ;
        RECT  5.770 3.545 6.000 4.365 ;
        RECT  5.635 0.955 5.865 2.965 ;
        RECT  5.420 4.135 5.770 4.365 ;
        RECT  5.310 0.955 5.635 1.240 ;
        RECT  5.335 2.735 5.635 2.965 ;
        RECT  5.175 1.770 5.405 2.225 ;
        RECT  5.105 2.735 5.335 3.820 ;
        RECT  4.970 0.900 5.310 1.240 ;
        RECT  4.710 1.995 5.175 2.225 ;
        RECT  4.710 3.280 4.785 3.645 ;
        RECT  4.510 1.455 4.710 3.645 ;
        RECT  4.495 1.400 4.510 3.645 ;
        RECT  4.330 0.695 4.505 0.925 ;
        RECT  4.480 1.400 4.495 3.535 ;
        RECT  4.170 1.400 4.480 1.740 ;
        RECT  3.835 3.250 4.480 3.535 ;
        RECT  4.100 0.695 4.330 1.095 ;
        RECT  4.075 3.945 4.305 4.320 ;
        RECT  2.860 0.865 4.100 1.095 ;
        RECT  3.255 3.945 4.075 4.175 ;
        RECT  3.025 3.615 3.255 4.175 ;
        RECT  2.295 3.615 3.025 3.845 ;
        RECT  2.630 0.865 2.860 1.585 ;
        RECT  2.490 1.355 2.630 1.585 ;
        RECT  1.455 4.145 2.535 4.375 ;
        RECT  2.260 1.355 2.490 1.960 ;
        RECT  2.065 3.300 2.295 3.845 ;
        RECT  2.005 0.675 2.185 0.905 ;
        RECT  1.955 3.300 2.065 3.640 ;
        RECT  1.775 0.675 2.005 1.625 ;
        RECT  1.570 1.395 1.775 1.625 ;
        RECT  1.340 1.395 1.570 2.490 ;
        RECT  1.225 3.945 1.455 4.375 ;
        RECT  1.230 2.150 1.340 2.490 ;
        RECT  0.455 2.255 1.230 2.485 ;
        RECT  0.455 3.945 1.225 4.175 ;
        RECT  0.225 2.255 0.455 4.175 ;
    END
END SDFFSRX1

MACRO SDFFSHQXL
    CLASS CORE ;
    FOREIGN SDFFSHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 2.190 13.945 2.530 ;
        RECT  13.605 2.190 13.645 2.635 ;
        RECT  13.495 2.220 13.605 2.635 ;
        RECT  13.265 2.220 13.495 4.175 ;
        RECT  8.055 3.945 13.265 4.175 ;
        RECT  7.825 2.660 8.055 4.175 ;
        RECT  7.705 2.660 7.825 2.945 ;
        RECT  7.475 2.405 7.705 2.945 ;
        RECT  6.805 2.555 7.475 2.945 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.825 3.260 2.245 ;
        RECT  2.595 2.015 2.855 2.245 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.325 2.480 3.555 3.280 ;
        RECT  3.085 2.940 3.325 3.280 ;
        RECT  2.425 3.050 3.085 3.280 ;
        RECT  2.325 2.965 2.425 3.280 ;
        RECT  2.095 2.580 2.325 3.280 ;
        RECT  1.540 2.580 2.095 2.810 ;
        RECT  1.310 2.430 1.540 2.810 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.395 1.120 15.625 3.005 ;
        RECT  15.135 1.120 15.395 1.460 ;
        RECT  15.320 2.635 15.395 3.005 ;
        RECT  14.465 2.775 15.320 3.005 ;
        RECT  14.235 2.775 14.465 3.460 ;
        RECT  14.125 3.120 14.235 3.460 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.475 4.420 1.955 ;
        RECT  4.175 1.475 4.405 2.075 ;
        RECT  3.975 1.475 4.175 2.035 ;
        RECT  3.890 1.475 3.975 1.955 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.515 0.885 0.525 1.225 ;
        RECT  0.130 0.680 0.515 1.225 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.195 -0.400 15.840 0.400 ;
        RECT  13.855 -0.400 14.195 1.430 ;
        RECT  12.490 -0.400 13.855 0.400 ;
        RECT  12.150 -0.400 12.490 0.575 ;
        RECT  9.505 -0.400 12.150 0.400 ;
        RECT  9.275 -0.400 9.505 1.495 ;
        RECT  6.680 -0.400 9.275 0.400 ;
        RECT  6.340 -0.400 6.680 0.845 ;
        RECT  3.180 -0.400 6.340 0.400 ;
        RECT  2.840 -0.400 3.180 0.575 ;
        RECT  1.120 -0.400 2.840 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.185 4.640 15.840 5.440 ;
        RECT  14.845 3.320 15.185 5.440 ;
        RECT  13.855 4.640 14.845 5.440 ;
        RECT  13.515 4.465 13.855 5.440 ;
        RECT  12.475 4.640 13.515 5.440 ;
        RECT  12.135 4.465 12.475 5.440 ;
        RECT  9.300 4.640 12.135 5.440 ;
        RECT  8.935 4.465 9.300 5.440 ;
        RECT  7.590 4.640 8.935 5.440 ;
        RECT  6.650 4.140 7.590 5.440 ;
        RECT  3.400 4.640 6.650 5.440 ;
        RECT  3.060 4.465 3.400 5.440 ;
        RECT  1.100 4.640 3.060 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.080 2.165 15.085 2.450 ;
        RECT  14.855 1.725 15.080 2.450 ;
        RECT  14.850 1.725 14.855 2.395 ;
        RECT  13.245 1.725 14.850 1.955 ;
        RECT  13.130 0.805 13.245 1.955 ;
        RECT  13.015 0.695 13.130 1.955 ;
        RECT  12.775 0.695 13.015 1.040 ;
        RECT  12.780 2.640 12.985 3.150 ;
        RECT  12.755 1.290 12.780 3.150 ;
        RECT  12.200 0.810 12.775 1.040 ;
        RECT  12.550 1.290 12.755 2.870 ;
        RECT  11.890 2.640 12.550 2.870 ;
        RECT  11.970 0.810 12.200 2.265 ;
        RECT  11.125 0.810 11.970 1.040 ;
        RECT  11.430 2.035 11.970 2.265 ;
        RECT  11.660 2.640 11.890 3.000 ;
        RECT  11.200 1.430 11.540 1.770 ;
        RECT  9.365 3.440 11.505 3.670 ;
        RECT  11.200 2.035 11.430 3.190 ;
        RECT  10.970 1.540 11.200 1.770 ;
        RECT  10.560 2.960 11.200 3.190 ;
        RECT  10.785 0.755 11.125 1.095 ;
        RECT  10.740 1.540 10.970 2.445 ;
        RECT  10.350 2.215 10.740 2.445 ;
        RECT  10.255 1.105 10.365 1.445 ;
        RECT  10.120 2.215 10.350 2.580 ;
        RECT  10.025 1.105 10.255 1.965 ;
        RECT  9.875 2.960 10.050 3.190 ;
        RECT  9.875 1.735 10.025 1.965 ;
        RECT  9.645 1.735 9.875 3.190 ;
        RECT  9.135 1.870 9.365 3.670 ;
        RECT  9.035 1.870 9.135 2.100 ;
        RECT  9.015 3.395 9.135 3.670 ;
        RECT  8.805 1.350 9.035 2.100 ;
        RECT  8.625 3.395 9.015 3.625 ;
        RECT  8.575 2.330 8.900 2.670 ;
        RECT  8.705 1.350 8.805 1.580 ;
        RECT  8.475 0.675 8.705 1.580 ;
        RECT  8.285 3.340 8.625 3.680 ;
        RECT  8.560 1.810 8.575 2.670 ;
        RECT  8.345 1.810 8.560 2.615 ;
        RECT  8.140 0.675 8.475 0.905 ;
        RECT  8.190 1.810 8.345 2.040 ;
        RECT  7.960 1.335 8.190 2.040 ;
        RECT  7.600 1.335 7.960 1.995 ;
        RECT  7.265 0.775 7.705 1.005 ;
        RECT  6.575 1.765 7.600 1.995 ;
        RECT  6.575 3.395 7.300 3.625 ;
        RECT  7.035 0.775 7.265 1.365 ;
        RECT  5.630 1.135 7.035 1.365 ;
        RECT  6.345 1.765 6.575 3.625 ;
        RECT  5.955 1.885 6.345 2.115 ;
        RECT  5.885 2.360 6.115 3.635 ;
        RECT  5.625 2.360 5.885 2.590 ;
        RECT  5.415 3.405 5.885 3.635 ;
        RECT  4.980 2.825 5.655 3.055 ;
        RECT  5.625 1.015 5.630 1.365 ;
        RECT  5.395 1.015 5.625 2.590 ;
        RECT  5.075 3.405 5.415 3.745 ;
        RECT  4.975 1.015 5.395 1.245 ;
        RECT  4.750 1.535 4.980 3.055 ;
        RECT  4.120 2.825 4.750 3.055 ;
        RECT  4.360 3.550 4.590 4.230 ;
        RECT  4.165 0.720 4.505 1.060 ;
        RECT  1.650 4.000 4.360 4.230 ;
        RECT  1.765 0.815 4.165 1.045 ;
        RECT  3.890 2.825 4.120 3.765 ;
        RECT  0.520 3.535 3.890 3.765 ;
        RECT  2.025 1.335 3.540 1.565 ;
        RECT  2.025 1.900 2.210 2.340 ;
        RECT  1.980 1.335 2.025 2.340 ;
        RECT  1.795 1.335 1.980 2.200 ;
        RECT  0.985 3.075 1.865 3.305 ;
        RECT  1.680 1.455 1.795 2.200 ;
        RECT  1.535 0.640 1.765 1.045 ;
        RECT  0.985 1.970 1.680 2.200 ;
        RECT  0.755 1.970 0.985 3.305 ;
        RECT  0.370 3.150 0.520 3.765 ;
        RECT  0.370 1.455 0.465 1.915 ;
        RECT  0.290 1.455 0.370 3.765 ;
        RECT  0.235 1.455 0.290 3.490 ;
        RECT  0.180 1.685 0.235 3.490 ;
        RECT  0.140 1.685 0.180 3.390 ;
    END
END SDFFSHQXL

MACRO SDFFSHQX4
    CLASS CORE ;
    FOREIGN SDFFSHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSHQXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.355 2.250 19.580 2.480 ;
        RECT  19.020 2.250 19.355 2.565 ;
        RECT  17.695 2.335 19.020 2.565 ;
        RECT  17.650 2.255 17.695 2.565 ;
        RECT  17.420 2.255 17.650 4.235 ;
        RECT  17.280 2.255 17.420 2.485 ;
        RECT  17.300 3.755 17.420 4.235 ;
        RECT  12.685 4.005 17.300 4.235 ;
        RECT  12.455 3.530 12.685 4.235 ;
        RECT  8.285 3.530 12.455 3.760 ;
        RECT  8.285 2.965 8.365 3.195 ;
        RECT  8.055 2.900 8.285 3.760 ;
        RECT  7.070 2.900 8.055 3.130 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.500 3.155 2.840 ;
        RECT  2.855 1.350 3.085 2.840 ;
        RECT  2.720 1.350 2.855 1.580 ;
        RECT  2.815 2.500 2.855 2.840 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.720 2.405 1.765 2.715 ;
        RECT  1.260 2.380 1.720 2.810 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.920 0.800 20.940 1.285 ;
        RECT  20.690 0.800 20.920 3.185 ;
        RECT  20.600 0.800 20.690 1.495 ;
        RECT  20.320 2.955 20.690 3.185 ;
        RECT  18.380 1.265 20.600 1.495 ;
        RECT  19.940 2.940 20.320 4.340 ;
        RECT  19.720 2.985 19.940 4.030 ;
        RECT  19.585 2.985 19.720 3.220 ;
        RECT  18.695 2.985 19.585 3.215 ;
        RECT  18.540 2.985 18.695 3.220 ;
        RECT  18.200 2.985 18.540 3.925 ;
        RECT  18.145 1.055 18.380 1.495 ;
        RECT  18.040 1.055 18.145 1.395 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.380 4.480 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 1.755 1.250 2.140 ;
        RECT  0.695 1.755 0.925 2.330 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.660 -0.400 21.120 0.400 ;
        RECT  19.320 -0.400 19.660 0.955 ;
        RECT  15.740 -0.400 19.320 0.400 ;
        RECT  15.400 -0.400 15.740 0.575 ;
        RECT  11.460 -0.400 15.400 0.400 ;
        RECT  11.120 -0.400 11.460 1.280 ;
        RECT  10.015 -0.400 11.120 0.400 ;
        RECT  9.675 -0.400 10.015 1.395 ;
        RECT  6.725 -0.400 9.675 0.400 ;
        RECT  6.385 -0.400 6.725 1.040 ;
        RECT  3.440 -0.400 6.385 0.400 ;
        RECT  3.100 -0.400 3.440 0.575 ;
        RECT  1.295 -0.400 3.100 0.400 ;
        RECT  0.955 -0.400 1.295 0.575 ;
        RECT  0.000 -0.400 0.955 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.855 4.640 21.120 5.440 ;
        RECT  20.625 3.480 20.855 5.440 ;
        RECT  19.300 4.640 20.625 5.440 ;
        RECT  18.960 3.480 19.300 5.440 ;
        RECT  17.740 4.640 18.960 5.440 ;
        RECT  17.400 4.465 17.740 5.440 ;
        RECT  16.270 4.640 17.400 5.440 ;
        RECT  15.930 4.465 16.270 5.440 ;
        RECT  11.590 4.640 15.930 5.440 ;
        RECT  11.250 4.465 11.590 5.440 ;
        RECT  10.065 4.640 11.250 5.440 ;
        RECT  9.725 4.465 10.065 5.440 ;
        RECT  8.600 4.640 9.725 5.440 ;
        RECT  8.260 4.465 8.600 5.440 ;
        RECT  7.080 4.640 8.260 5.440 ;
        RECT  6.740 4.465 7.080 5.440 ;
        RECT  3.805 4.640 6.740 5.440 ;
        RECT  3.465 4.155 3.805 5.440 ;
        RECT  1.300 4.640 3.465 5.440 ;
        RECT  0.960 4.465 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.350 2.205 20.460 2.545 ;
        RECT  20.120 1.780 20.350 2.545 ;
        RECT  18.720 1.780 20.120 2.010 ;
        RECT  18.320 1.780 18.720 2.065 ;
        RECT  17.655 1.780 18.320 2.010 ;
        RECT  17.425 0.865 17.655 2.010 ;
        RECT  14.845 0.865 17.425 1.095 ;
        RECT  16.950 3.000 17.060 3.340 ;
        RECT  16.720 1.545 16.950 3.340 ;
        RECT  15.900 1.545 16.720 1.775 ;
        RECT  16.345 2.250 16.455 2.590 ;
        RECT  16.115 2.250 16.345 3.775 ;
        RECT  14.845 3.545 16.115 3.775 ;
        RECT  15.560 1.410 15.900 1.775 ;
        RECT  15.525 1.540 15.560 1.775 ;
        RECT  15.240 1.540 15.525 2.345 ;
        RECT  15.185 2.005 15.240 2.345 ;
        RECT  14.615 0.865 14.845 3.775 ;
        RECT  14.340 0.865 14.615 1.095 ;
        RECT  13.060 3.545 14.615 3.775 ;
        RECT  14.230 0.865 14.340 1.410 ;
        RECT  14.000 0.725 14.230 1.410 ;
        RECT  13.520 3.070 14.160 3.300 ;
        RECT  12.900 0.725 14.000 0.955 ;
        RECT  13.520 1.200 13.620 1.540 ;
        RECT  13.290 1.200 13.520 3.300 ;
        RECT  13.280 1.200 13.290 1.745 ;
        RECT  12.270 3.070 13.290 3.300 ;
        RECT  12.180 1.515 13.280 1.745 ;
        RECT  12.670 0.725 12.900 1.275 ;
        RECT  12.560 0.935 12.670 1.275 ;
        RECT  9.945 1.975 12.665 2.205 ;
        RECT  12.040 2.985 12.270 3.300 ;
        RECT  11.840 1.100 12.180 1.745 ;
        RECT  11.895 3.995 12.125 4.405 ;
        RECT  10.825 2.985 12.040 3.215 ;
        RECT  6.135 3.995 11.895 4.225 ;
        RECT  10.740 1.515 11.840 1.745 ;
        RECT  10.485 2.875 10.825 3.215 ;
        RECT  10.455 1.110 10.740 1.745 ;
        RECT  10.400 1.110 10.455 1.450 ;
        RECT  9.715 1.805 9.945 3.155 ;
        RECT  9.225 1.805 9.715 2.035 ;
        RECT  9.445 2.870 9.715 3.155 ;
        RECT  8.275 2.295 9.470 2.525 ;
        RECT  9.105 2.870 9.445 3.210 ;
        RECT  8.995 0.775 9.225 2.035 ;
        RECT  7.490 0.775 8.995 1.005 ;
        RECT  8.205 1.300 8.275 2.665 ;
        RECT  8.045 1.245 8.205 2.665 ;
        RECT  7.865 1.245 8.045 1.585 ;
        RECT  6.505 2.435 8.045 2.665 ;
        RECT  5.840 1.975 7.815 2.205 ;
        RECT  7.555 3.365 7.785 3.760 ;
        RECT  6.505 3.365 7.555 3.595 ;
        RECT  7.260 0.775 7.490 1.705 ;
        RECT  6.125 1.475 7.260 1.705 ;
        RECT  6.275 2.435 6.505 3.595 ;
        RECT  5.850 3.995 6.135 4.235 ;
        RECT  5.895 0.635 6.125 1.705 ;
        RECT  5.715 0.635 5.895 0.865 ;
        RECT  5.375 4.005 5.850 4.235 ;
        RECT  5.610 1.975 5.840 3.715 ;
        RECT  5.485 1.975 5.610 2.205 ;
        RECT  5.255 0.830 5.485 2.205 ;
        RECT  5.145 3.075 5.375 4.235 ;
        RECT  5.140 0.830 5.255 1.060 ;
        RECT  5.015 3.075 5.145 3.305 ;
        RECT  4.785 1.455 5.015 3.305 ;
        RECT  4.625 3.595 4.855 4.050 ;
        RECT  2.765 3.075 4.785 3.305 ;
        RECT  2.040 0.815 4.760 1.045 ;
        RECT  3.230 3.595 4.625 3.825 ;
        RECT  3.000 3.595 3.230 4.295 ;
        RECT  1.940 4.065 3.000 4.295 ;
        RECT  2.535 3.075 2.765 3.835 ;
        RECT  0.530 3.605 2.535 3.835 ;
        RECT  2.300 2.070 2.415 2.410 ;
        RECT  2.070 1.570 2.300 3.315 ;
        RECT  2.055 1.570 2.070 1.800 ;
        RECT  1.620 3.085 2.070 3.315 ;
        RECT  1.715 1.460 2.055 1.800 ;
        RECT  1.755 0.650 2.040 1.045 ;
        RECT  1.700 0.650 1.755 0.990 ;
        RECT  0.420 1.180 0.530 1.520 ;
        RECT  0.420 3.000 0.530 3.940 ;
        RECT  0.190 1.180 0.420 3.940 ;
    END
END SDFFSHQX4

MACRO SDFFSHQX2
    CLASS CORE ;
    FOREIGN SDFFSHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSHQXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.545 2.110 17.775 3.755 ;
        RECT  15.355 3.525 17.545 3.755 ;
        RECT  15.355 2.175 15.420 2.515 ;
        RECT  15.125 2.175 15.355 3.755 ;
        RECT  15.080 2.175 15.125 2.515 ;
        RECT  15.050 3.525 15.125 3.755 ;
        RECT  14.820 3.525 15.050 4.305 ;
        RECT  11.000 4.075 14.820 4.305 ;
        RECT  10.770 3.655 11.000 4.305 ;
        RECT  10.700 3.655 10.770 4.085 ;
        RECT  9.760 3.655 10.700 3.885 ;
        RECT  9.570 3.655 9.760 4.085 ;
        RECT  9.340 3.655 9.570 4.365 ;
        RECT  7.785 4.135 9.340 4.365 ;
        RECT  7.705 2.455 7.785 4.365 ;
        RECT  7.555 2.405 7.705 4.365 ;
        RECT  6.755 2.405 7.555 2.685 ;
        RECT  6.470 2.405 6.755 2.780 ;
        RECT  6.415 2.440 6.470 2.780 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.615 2.300 3.135 2.760 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 2.035 1.610 2.375 ;
        RECT  1.270 1.865 1.305 2.375 ;
        RECT  1.105 1.865 1.270 2.320 ;
        RECT  1.075 1.845 1.105 2.320 ;
        RECT  0.875 1.845 1.075 2.095 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.055 1.290 17.285 3.080 ;
        RECT  16.945 1.290 17.055 1.540 ;
        RECT  16.715 2.850 17.055 3.080 ;
        RECT  16.850 1.290 16.945 1.520 ;
        RECT  16.510 1.180 16.850 1.520 ;
        RECT  16.380 2.850 16.715 3.190 ;
        RECT  16.055 2.850 16.380 3.195 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 1.825 3.985 2.340 ;
        RECT  3.515 1.845 3.565 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 3.805 0.675 4.235 ;
        RECT  0.215 3.805 0.475 4.315 ;
        RECT  0.190 3.805 0.215 4.235 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.130 -0.400 18.480 0.400 ;
        RECT  17.790 -0.400 18.130 1.510 ;
        RECT  14.445 -0.400 17.790 0.400 ;
        RECT  14.105 -0.400 14.445 0.575 ;
        RECT  10.925 -0.400 14.105 0.400 ;
        RECT  10.585 -0.400 10.925 1.335 ;
        RECT  9.430 -0.400 10.585 0.400 ;
        RECT  9.200 -0.400 9.430 1.370 ;
        RECT  6.505 -0.400 9.200 0.400 ;
        RECT  6.165 -0.400 6.505 0.960 ;
        RECT  3.140 -0.400 6.165 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.080 -0.400 2.800 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.155 4.640 18.480 5.440 ;
        RECT  16.815 4.085 17.155 5.440 ;
        RECT  15.655 4.640 16.815 5.440 ;
        RECT  15.315 4.035 15.655 5.440 ;
        RECT  10.390 4.640 15.315 5.440 ;
        RECT  10.050 4.120 10.390 5.440 ;
        RECT  7.325 4.640 10.050 5.440 ;
        RECT  6.515 4.140 7.325 5.440 ;
        RECT  3.375 4.640 6.515 5.440 ;
        RECT  3.035 4.140 3.375 5.440 ;
        RECT  1.090 4.640 3.035 5.440 ;
        RECT  0.750 4.465 1.090 5.440 ;
        RECT  0.000 4.640 0.750 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.890 2.095 16.705 2.325 ;
        RECT  15.660 0.865 15.890 2.325 ;
        RECT  13.115 0.865 15.660 1.095 ;
        RECT  14.410 2.125 14.590 3.745 ;
        RECT  14.360 2.125 14.410 3.800 ;
        RECT  14.285 2.125 14.360 2.355 ;
        RECT  14.070 3.460 14.360 3.800 ;
        RECT  14.285 1.460 14.340 1.800 ;
        RECT  14.055 1.460 14.285 2.355 ;
        RECT  13.785 2.760 14.125 3.100 ;
        RECT  14.000 1.460 14.055 1.800 ;
        RECT  14.040 2.060 14.055 2.355 ;
        RECT  13.700 2.060 14.040 2.400 ;
        RECT  13.115 2.815 13.785 3.045 ;
        RECT  12.955 0.865 13.115 3.845 ;
        RECT  12.885 0.795 12.955 3.845 ;
        RECT  12.725 0.795 12.885 1.600 ;
        RECT  11.530 3.615 12.885 3.845 ;
        RECT  11.625 0.795 12.725 1.025 ;
        RECT  12.395 3.135 12.650 3.365 ;
        RECT  12.345 1.595 12.395 3.365 ;
        RECT  12.165 1.280 12.345 3.365 ;
        RECT  12.005 1.280 12.165 1.825 ;
        RECT  11.150 3.135 12.165 3.365 ;
        RECT  10.205 1.595 12.005 1.825 ;
        RECT  9.105 2.055 11.925 2.285 ;
        RECT  11.395 0.795 11.625 1.365 ;
        RECT  11.285 1.025 11.395 1.365 ;
        RECT  10.810 3.080 11.150 3.420 ;
        RECT  9.675 3.135 10.810 3.365 ;
        RECT  9.975 1.115 10.205 1.825 ;
        RECT  9.865 1.115 9.975 1.455 ;
        RECT  9.335 3.080 9.675 3.420 ;
        RECT  8.875 1.750 9.105 3.845 ;
        RECT  8.730 1.750 8.875 1.980 ;
        RECT  8.695 3.505 8.875 3.845 ;
        RECT  8.630 1.410 8.730 1.980 ;
        RECT  8.485 3.560 8.695 3.845 ;
        RECT  8.500 0.675 8.630 1.980 ;
        RECT  8.390 2.240 8.620 2.875 ;
        RECT  8.400 0.675 8.500 1.640 ;
        RECT  8.145 3.560 8.485 3.900 ;
        RECT  7.985 0.675 8.400 0.905 ;
        RECT  8.260 2.240 8.390 2.470 ;
        RECT  8.030 1.875 8.260 2.470 ;
        RECT  7.885 1.875 8.030 2.105 ;
        RECT  7.655 1.415 7.885 2.105 ;
        RECT  7.545 1.415 7.655 1.885 ;
        RECT  7.305 0.720 7.645 1.060 ;
        RECT  6.025 1.655 7.545 1.885 ;
        RECT  7.185 0.830 7.305 1.060 ;
        RECT  6.955 0.830 7.185 1.420 ;
        RECT  6.820 3.270 7.160 3.610 ;
        RECT  5.220 1.190 6.955 1.420 ;
        RECT  6.025 3.325 6.820 3.555 ;
        RECT  6.025 2.170 6.080 2.510 ;
        RECT  5.795 1.655 6.025 3.555 ;
        RECT  5.740 2.170 5.795 2.510 ;
        RECT  5.275 3.905 5.615 4.245 ;
        RECT  4.760 3.960 5.275 4.190 ;
        RECT  4.990 1.190 5.220 3.570 ;
        RECT  4.780 1.355 4.990 1.585 ;
        RECT  4.650 3.075 4.760 4.190 ;
        RECT  4.650 1.855 4.705 2.195 ;
        RECT  4.530 1.855 4.650 4.190 ;
        RECT  4.425 0.655 4.560 0.885 ;
        RECT  4.420 1.855 4.530 3.305 ;
        RECT  4.195 0.655 4.425 1.095 ;
        RECT  4.365 1.855 4.420 2.195 ;
        RECT  2.245 3.075 4.420 3.305 ;
        RECT  4.070 3.595 4.300 4.110 ;
        RECT  1.780 0.865 4.195 1.095 ;
        RECT  2.750 3.595 4.070 3.825 ;
        RECT  2.235 1.325 3.470 1.555 ;
        RECT  2.520 3.595 2.750 4.295 ;
        RECT  1.670 4.065 2.520 4.295 ;
        RECT  2.015 3.075 2.245 3.835 ;
        RECT  2.005 1.325 2.235 2.845 ;
        RECT  1.320 3.605 2.015 3.835 ;
        RECT  1.985 1.325 2.005 1.780 ;
        RECT  1.785 2.615 2.005 2.845 ;
        RECT  1.540 1.440 1.985 1.780 ;
        RECT  1.555 2.615 1.785 3.270 ;
        RECT  1.550 0.630 1.780 1.095 ;
        RECT  1.440 0.630 1.550 0.970 ;
        RECT  1.090 3.245 1.320 3.835 ;
        RECT  0.520 3.245 1.090 3.475 ;
        RECT  0.375 1.355 0.520 1.695 ;
        RECT  0.375 3.135 0.520 3.475 ;
        RECT  0.180 1.355 0.375 3.475 ;
        RECT  0.145 1.465 0.180 3.420 ;
    END
END SDFFSHQX2

MACRO SDFFSHQX1
    CLASS CORE ;
    FOREIGN SDFFSHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSHQXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.075 1.845 14.305 2.100 ;
        RECT  13.945 1.870 14.075 2.100 ;
        RECT  13.715 1.870 13.945 2.450 ;
        RECT  13.605 2.110 13.715 2.450 ;
        RECT  13.495 2.220 13.605 2.450 ;
        RECT  13.265 2.220 13.495 4.175 ;
        RECT  8.055 3.945 13.265 4.175 ;
        RECT  7.825 2.660 8.055 4.175 ;
        RECT  7.705 2.660 7.825 2.945 ;
        RECT  7.475 2.405 7.705 2.945 ;
        RECT  6.805 2.555 7.475 2.945 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.055 1.445 3.085 2.775 ;
        RECT  2.990 1.445 3.055 2.830 ;
        RECT  2.855 1.390 2.990 2.830 ;
        RECT  2.780 1.390 2.855 1.845 ;
        RECT  2.715 2.490 2.855 2.830 ;
        RECT  2.650 1.390 2.780 1.730 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 2.265 1.870 2.810 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.395 0.855 15.625 3.005 ;
        RECT  15.320 0.855 15.395 1.290 ;
        RECT  15.320 2.635 15.395 3.005 ;
        RECT  15.190 0.855 15.320 1.220 ;
        RECT  14.465 2.775 15.320 3.005 ;
        RECT  14.235 2.775 14.465 3.440 ;
        RECT  14.125 3.100 14.235 3.440 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.890 1.770 4.420 2.250 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 1.845 1.105 2.075 ;
        RECT  1.015 1.845 1.030 2.375 ;
        RECT  0.835 1.845 1.015 2.380 ;
        RECT  0.785 1.845 0.835 2.510 ;
        RECT  0.605 2.145 0.785 2.510 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.155 -0.400 15.840 0.400 ;
        RECT  13.815 -0.400 14.155 0.575 ;
        RECT  12.490 -0.400 13.815 0.400 ;
        RECT  12.150 -0.400 12.490 0.575 ;
        RECT  9.505 -0.400 12.150 0.400 ;
        RECT  9.275 -0.400 9.505 1.280 ;
        RECT  6.680 -0.400 9.275 0.400 ;
        RECT  6.340 -0.400 6.680 0.845 ;
        RECT  3.150 -0.400 6.340 0.400 ;
        RECT  2.810 -0.400 3.150 0.575 ;
        RECT  1.080 -0.400 2.810 0.400 ;
        RECT  0.740 -0.400 1.080 0.930 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.185 4.640 15.840 5.440 ;
        RECT  14.845 3.320 15.185 5.440 ;
        RECT  13.880 4.640 14.845 5.440 ;
        RECT  13.540 4.465 13.880 5.440 ;
        RECT  12.475 4.640 13.540 5.440 ;
        RECT  12.135 4.465 12.475 5.440 ;
        RECT  9.300 4.640 12.135 5.440 ;
        RECT  8.935 4.465 9.300 5.440 ;
        RECT  7.590 4.640 8.935 5.440 ;
        RECT  6.650 4.140 7.590 5.440 ;
        RECT  3.720 4.640 6.650 5.440 ;
        RECT  3.490 4.145 3.720 5.440 ;
        RECT  1.100 4.640 3.490 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.950 2.110 15.060 2.450 ;
        RECT  14.720 1.285 14.950 2.450 ;
        RECT  13.245 1.285 14.720 1.515 ;
        RECT  13.130 0.805 13.245 1.515 ;
        RECT  13.015 0.695 13.130 1.515 ;
        RECT  12.795 2.640 13.025 3.150 ;
        RECT  12.775 0.695 13.015 1.035 ;
        RECT  12.780 2.640 12.795 2.870 ;
        RECT  12.550 1.320 12.780 2.870 ;
        RECT  12.020 0.805 12.775 1.035 ;
        RECT  11.945 2.640 12.550 2.870 ;
        RECT  11.790 0.805 12.020 2.265 ;
        RECT  11.605 2.640 11.945 2.980 ;
        RECT  11.305 0.805 11.790 1.035 ;
        RECT  11.210 2.035 11.790 2.265 ;
        RECT  10.740 1.450 11.540 1.680 ;
        RECT  9.365 3.440 11.505 3.670 ;
        RECT  11.070 0.805 11.305 1.220 ;
        RECT  10.980 2.035 11.210 3.190 ;
        RECT  10.665 0.990 11.070 1.220 ;
        RECT  10.560 2.960 10.980 3.190 ;
        RECT  10.510 1.450 10.740 2.445 ;
        RECT  10.350 2.215 10.510 2.445 ;
        RECT  10.120 2.215 10.350 2.580 ;
        RECT  10.170 1.080 10.280 1.420 ;
        RECT  9.940 1.080 10.170 1.835 ;
        RECT  9.875 2.960 10.095 3.190 ;
        RECT  9.875 1.605 9.940 1.835 ;
        RECT  9.645 1.605 9.875 3.190 ;
        RECT  9.135 1.595 9.365 3.670 ;
        RECT  9.035 1.595 9.135 1.825 ;
        RECT  9.015 3.375 9.135 3.670 ;
        RECT  8.805 1.350 9.035 1.825 ;
        RECT  8.625 3.375 9.015 3.660 ;
        RECT  8.575 2.355 8.900 2.585 ;
        RECT  8.760 1.350 8.805 1.580 ;
        RECT  8.650 1.240 8.760 1.580 ;
        RECT  8.480 0.685 8.650 1.580 ;
        RECT  8.285 3.320 8.625 3.660 ;
        RECT  8.345 1.810 8.575 2.585 ;
        RECT  8.420 0.630 8.480 1.580 ;
        RECT  8.140 0.630 8.420 0.970 ;
        RECT  8.075 1.810 8.345 2.040 ;
        RECT  7.845 1.335 8.075 2.040 ;
        RECT  7.695 1.335 7.845 1.995 ;
        RECT  7.365 0.720 7.705 1.060 ;
        RECT  6.575 1.765 7.695 1.995 ;
        RECT  7.265 0.830 7.365 1.060 ;
        RECT  6.960 3.340 7.300 3.680 ;
        RECT  7.035 0.830 7.265 1.365 ;
        RECT  5.630 1.135 7.035 1.365 ;
        RECT  6.575 3.340 6.960 3.570 ;
        RECT  6.345 1.765 6.575 3.570 ;
        RECT  5.955 1.790 6.345 2.130 ;
        RECT  5.885 2.365 6.115 3.850 ;
        RECT  5.625 2.365 5.885 2.595 ;
        RECT  5.375 3.620 5.885 3.850 ;
        RECT  5.315 2.940 5.655 3.280 ;
        RECT  5.625 0.855 5.630 1.365 ;
        RECT  5.395 0.855 5.625 2.595 ;
        RECT  5.315 0.855 5.395 1.140 ;
        RECT  5.035 3.620 5.375 3.960 ;
        RECT  4.975 0.800 5.315 1.140 ;
        RECT  5.000 2.940 5.315 3.170 ;
        RECT  5.000 1.840 5.055 2.180 ;
        RECT  4.770 1.840 5.000 3.170 ;
        RECT  4.715 1.840 4.770 2.180 ;
        RECT  3.690 2.525 4.770 2.755 ;
        RECT  4.235 3.465 4.575 3.805 ;
        RECT  4.460 1.080 4.510 1.420 ;
        RECT  4.170 0.865 4.460 1.420 ;
        RECT  3.255 3.575 4.235 3.805 ;
        RECT  1.725 0.865 4.170 1.095 ;
        RECT  3.460 2.525 3.690 3.305 ;
        RECT  2.790 3.075 3.460 3.305 ;
        RECT  3.025 3.575 3.255 4.305 ;
        RECT  1.650 4.075 3.025 4.305 ;
        RECT  2.560 3.075 2.790 3.845 ;
        RECT  0.520 3.615 2.560 3.845 ;
        RECT  2.100 1.635 2.330 3.315 ;
        RECT  2.020 1.635 2.100 1.865 ;
        RECT  1.525 3.085 2.100 3.315 ;
        RECT  1.735 1.455 2.020 1.865 ;
        RECT  1.680 1.455 1.735 1.795 ;
        RECT  1.495 0.640 1.725 1.095 ;
        RECT  0.370 1.390 0.520 1.730 ;
        RECT  0.370 3.120 0.520 3.845 ;
        RECT  0.290 1.390 0.370 3.845 ;
        RECT  0.180 1.390 0.290 3.460 ;
        RECT  0.140 1.390 0.180 3.390 ;
    END
END SDFFSHQX1

MACRO SDFFSXL
    CLASS CORE ;
    FOREIGN SDFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.020 4.060 12.650 4.410 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.150 2.110 3.275 2.635 ;
        RECT  3.045 2.110 3.150 2.650 ;
        RECT  2.750 2.150 3.045 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.830 1.815 1.600 2.100 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.200 0.865 14.430 3.950 ;
        RECT  13.725 0.865 14.200 1.095 ;
        RECT  14.000 3.720 14.200 3.950 ;
        RECT  13.645 3.720 14.000 4.105 ;
        RECT  13.495 0.680 13.725 1.095 ;
        RECT  13.415 3.720 13.645 4.315 ;
        RECT  13.280 0.680 13.495 1.020 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.965 3.090 15.260 3.430 ;
        RECT  14.965 1.250 15.220 1.590 ;
        RECT  14.880 1.250 14.965 3.430 ;
        RECT  14.735 1.305 14.880 3.430 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 2.080 4.510 2.310 ;
        RECT  4.100 1.820 4.480 2.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.830 0.755 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.570 -0.400 15.840 0.400 ;
        RECT  14.230 -0.400 14.570 0.575 ;
        RECT  12.860 -0.400 14.230 0.400 ;
        RECT  12.520 -0.400 12.860 0.575 ;
        RECT  11.400 -0.400 12.520 0.400 ;
        RECT  11.060 -0.400 11.400 0.575 ;
        RECT  9.005 -0.400 11.060 0.400 ;
        RECT  8.775 -0.400 9.005 0.870 ;
        RECT  6.980 -0.400 8.775 0.400 ;
        RECT  6.640 -0.400 6.980 0.995 ;
        RECT  3.585 -0.400 6.640 0.400 ;
        RECT  3.245 -0.400 3.585 0.575 ;
        RECT  1.425 -0.400 3.245 0.400 ;
        RECT  1.085 -0.400 1.425 0.575 ;
        RECT  0.000 -0.400 1.085 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.745 4.640 15.840 5.440 ;
        RECT  14.345 4.465 14.745 5.440 ;
        RECT  13.110 4.640 14.345 5.440 ;
        RECT  13.110 2.920 13.280 3.260 ;
        RECT  12.940 2.920 13.110 5.440 ;
        RECT  12.880 2.975 12.940 5.440 ;
        RECT  11.790 4.640 12.880 5.440 ;
        RECT  11.450 4.140 11.790 5.440 ;
        RECT  9.280 4.640 11.450 5.440 ;
        RECT  8.940 4.140 9.280 5.440 ;
        RECT  7.965 4.640 8.940 5.440 ;
        RECT  7.735 4.140 7.965 5.440 ;
        RECT  6.620 4.640 7.735 5.440 ;
        RECT  6.280 4.465 6.620 5.440 ;
        RECT  3.485 4.640 6.280 5.440 ;
        RECT  3.255 4.100 3.485 5.440 ;
        RECT  1.080 4.640 3.255 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.945 1.545 13.970 2.940 ;
        RECT  13.740 1.545 13.945 3.260 ;
        RECT  13.660 1.545 13.740 1.775 ;
        RECT  13.715 2.710 13.740 3.260 ;
        RECT  13.320 1.435 13.660 1.775 ;
        RECT  12.520 2.025 13.355 2.255 ;
        RECT  12.325 1.895 12.520 3.380 ;
        RECT  12.290 1.515 12.325 3.380 ;
        RECT  12.095 1.515 12.290 2.125 ;
        RECT  12.180 3.040 12.290 3.380 ;
        RECT  11.700 1.515 12.095 1.745 ;
        RECT  10.545 2.435 12.040 2.665 ;
        RECT  11.360 1.405 11.700 1.745 ;
        RECT  11.050 1.405 11.360 1.635 ;
        RECT  10.815 1.160 11.050 1.635 ;
        RECT  10.710 1.160 10.815 1.500 ;
        RECT  10.545 3.290 10.600 3.630 ;
        RECT  10.475 1.875 10.545 3.630 ;
        RECT  10.315 1.495 10.475 3.630 ;
        RECT  10.250 1.495 10.315 2.105 ;
        RECT  10.260 3.290 10.315 3.630 ;
        RECT  10.245 1.440 10.250 2.105 ;
        RECT  9.910 1.440 10.245 1.780 ;
        RECT  9.890 4.020 10.230 4.360 ;
        RECT  9.775 2.015 9.940 2.355 ;
        RECT  9.740 4.020 9.890 4.250 ;
        RECT  9.680 2.015 9.775 3.145 ;
        RECT  9.510 3.670 9.740 4.250 ;
        RECT  9.450 1.245 9.680 3.145 ;
        RECT  6.245 3.670 9.510 3.900 ;
        RECT  8.545 1.245 9.450 1.475 ;
        RECT  8.725 2.915 9.450 3.145 ;
        RECT  8.875 2.165 9.215 2.505 ;
        RECT  8.265 2.220 8.875 2.450 ;
        RECT  8.495 2.915 8.725 3.420 ;
        RECT  8.315 0.725 8.545 1.475 ;
        RECT  8.035 0.725 8.315 0.955 ;
        RECT  8.085 2.220 8.265 3.415 ;
        RECT  8.035 1.450 8.085 3.415 ;
        RECT  7.805 0.635 8.035 0.955 ;
        RECT  7.855 1.450 8.035 2.450 ;
        RECT  6.470 3.185 8.035 3.415 ;
        RECT  7.310 0.635 7.805 0.865 ;
        RECT  7.230 2.445 7.570 2.785 ;
        RECT  6.930 2.445 7.230 2.675 ;
        RECT  6.700 2.180 6.930 2.675 ;
        RECT  5.690 2.180 6.700 2.410 ;
        RECT  6.240 2.640 6.470 3.415 ;
        RECT  6.015 3.670 6.245 4.085 ;
        RECT  6.120 2.640 6.240 2.870 ;
        RECT  5.685 3.855 6.015 4.085 ;
        RECT  5.690 0.680 5.745 1.020 ;
        RECT  5.460 0.680 5.690 3.125 ;
        RECT  5.400 3.855 5.685 4.405 ;
        RECT  5.405 0.680 5.460 1.020 ;
        RECT  5.445 2.895 5.460 3.125 ;
        RECT  5.215 2.895 5.445 3.520 ;
        RECT  4.985 4.175 5.400 4.405 ;
        RECT  5.170 1.400 5.225 1.740 ;
        RECT  4.985 1.400 5.170 2.430 ;
        RECT  4.940 1.400 4.985 4.405 ;
        RECT  4.605 0.760 4.945 1.100 ;
        RECT  4.885 1.400 4.940 1.740 ;
        RECT  4.755 2.200 4.940 4.405 ;
        RECT  3.945 4.175 4.755 4.405 ;
        RECT  2.640 0.870 4.605 1.100 ;
        RECT  4.405 3.715 4.525 3.945 ;
        RECT  4.175 3.035 4.405 3.945 ;
        RECT  2.425 3.035 4.175 3.265 ;
        RECT  3.715 3.630 3.945 4.405 ;
        RECT  2.415 1.405 3.865 1.635 ;
        RECT  3.020 3.630 3.715 3.860 ;
        RECT  2.790 3.630 3.020 4.365 ;
        RECT  1.685 4.135 2.790 4.365 ;
        RECT  2.410 0.695 2.640 1.100 ;
        RECT  2.415 2.465 2.470 2.805 ;
        RECT  2.380 3.035 2.425 3.845 ;
        RECT  2.225 1.405 2.415 2.805 ;
        RECT  1.885 0.695 2.410 0.925 ;
        RECT  2.195 3.035 2.380 3.900 ;
        RECT  2.185 1.350 2.225 2.805 ;
        RECT  2.040 3.560 2.195 3.900 ;
        RECT  1.885 1.350 2.185 1.690 ;
        RECT  2.130 2.465 2.185 2.805 ;
        RECT  1.825 2.575 2.130 2.805 ;
        RECT  1.595 2.575 1.825 3.160 ;
        RECT  1.455 3.650 1.685 4.365 ;
        RECT  1.215 3.650 1.455 3.880 ;
        RECT  0.985 2.350 1.215 3.880 ;
        RECT  0.410 2.350 0.985 2.580 ;
        RECT  0.180 3.540 0.985 3.880 ;
        RECT  0.410 1.190 0.520 1.530 ;
        RECT  0.180 1.190 0.410 2.580 ;
    END
END SDFFSXL

MACRO SDFFSX4
    CLASS CORE ;
    FOREIGN SDFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.170 4.040 7.780 4.410 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 2.050 3.250 2.635 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.820 1.765 2.500 ;
        RECT  1.410 2.075 1.460 2.500 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.000 1.360 19.020 1.700 ;
        RECT  19.000 2.740 19.020 3.080 ;
        RECT  18.660 1.260 19.000 3.080 ;
        RECT  18.620 1.260 18.660 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.830 1.820 20.980 3.220 ;
        RECT  20.600 1.470 20.830 3.220 ;
        RECT  20.300 1.470 20.600 1.700 ;
        RECT  19.960 2.740 20.600 3.080 ;
        RECT  19.960 1.360 20.300 1.700 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 1.840 4.405 2.365 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 2.380 1.180 2.660 ;
        RECT  0.720 1.835 0.950 2.660 ;
        RECT  0.610 1.835 0.720 2.175 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.940 -0.400 21.120 0.400 ;
        RECT  20.600 -0.400 20.940 0.950 ;
        RECT  19.660 -0.400 20.600 0.400 ;
        RECT  19.320 -0.400 19.660 0.950 ;
        RECT  18.340 -0.400 19.320 0.400 ;
        RECT  18.000 -0.400 18.340 0.575 ;
        RECT  16.990 -0.400 18.000 0.400 ;
        RECT  16.650 -0.400 16.990 1.100 ;
        RECT  14.390 -0.400 16.650 0.400 ;
        RECT  14.050 -0.400 14.390 0.575 ;
        RECT  12.400 -0.400 14.050 0.400 ;
        RECT  12.060 -0.400 12.400 1.320 ;
        RECT  9.840 -0.400 12.060 0.400 ;
        RECT  9.500 -0.400 9.840 1.320 ;
        RECT  6.920 -0.400 9.500 0.400 ;
        RECT  6.580 -0.400 6.920 1.280 ;
        RECT  3.400 -0.400 6.580 0.400 ;
        RECT  3.060 -0.400 3.400 0.575 ;
        RECT  1.180 -0.400 3.060 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.940 4.640 21.120 5.440 ;
        RECT  20.600 4.090 20.940 5.440 ;
        RECT  19.660 4.640 20.600 5.440 ;
        RECT  19.320 4.090 19.660 5.440 ;
        RECT  18.340 4.640 19.320 5.440 ;
        RECT  18.000 4.465 18.340 5.440 ;
        RECT  16.910 4.640 18.000 5.440 ;
        RECT  16.570 3.210 16.910 5.440 ;
        RECT  15.470 4.640 16.570 5.440 ;
        RECT  15.130 3.435 15.470 5.440 ;
        RECT  13.990 4.640 15.130 5.440 ;
        RECT  13.650 4.040 13.990 5.440 ;
        RECT  12.280 4.640 13.650 5.440 ;
        RECT  11.940 4.015 12.280 5.440 ;
        RECT  9.640 4.640 11.940 5.440 ;
        RECT  9.300 4.015 9.640 5.440 ;
        RECT  8.245 4.640 9.300 5.440 ;
        RECT  8.015 4.015 8.245 5.440 ;
        RECT  6.925 4.640 8.015 5.440 ;
        RECT  6.695 4.150 6.925 5.440 ;
        RECT  3.550 4.640 6.695 5.440 ;
        RECT  3.210 4.140 3.550 5.440 ;
        RECT  0.745 4.640 3.210 5.440 ;
        RECT  0.245 4.460 0.745 5.440 ;
        RECT  0.000 4.640 0.245 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.685 2.040 19.930 2.380 ;
        RECT  19.590 2.040 19.685 3.730 ;
        RECT  19.455 2.150 19.590 3.730 ;
        RECT  17.710 3.500 19.455 3.730 ;
        RECT  17.480 1.280 17.710 3.730 ;
        RECT  17.370 1.280 17.480 1.620 ;
        RECT  17.290 3.390 17.480 3.730 ;
        RECT  16.910 2.080 17.250 2.420 ;
        RECT  16.190 2.085 16.910 2.415 ;
        RECT  15.960 1.505 16.190 3.550 ;
        RECT  15.710 1.505 15.960 1.735 ;
        RECT  15.850 2.975 15.960 3.550 ;
        RECT  14.750 2.975 15.850 3.205 ;
        RECT  15.495 1.240 15.710 1.735 ;
        RECT  15.265 1.055 15.495 1.735 ;
        RECT  15.130 2.130 15.470 2.470 ;
        RECT  13.720 1.055 15.265 1.285 ;
        RECT  13.110 2.185 15.130 2.415 ;
        RECT  14.520 2.975 14.750 3.725 ;
        RECT  14.410 3.225 14.520 3.725 ;
        RECT  13.345 3.495 14.410 3.725 ;
        RECT  13.115 3.495 13.345 4.045 ;
        RECT  12.880 1.430 13.110 3.130 ;
        RECT  12.770 1.430 12.880 1.780 ;
        RECT  12.830 2.900 12.880 3.130 ;
        RECT  12.490 2.900 12.830 3.240 ;
        RECT  11.825 1.550 12.770 1.780 ;
        RECT  12.270 2.220 12.610 2.560 ;
        RECT  10.960 2.955 12.490 3.185 ;
        RECT  11.310 2.275 12.270 2.505 ;
        RECT  11.595 1.135 11.825 1.780 ;
        RECT  11.120 1.135 11.595 1.365 ;
        RECT  11.080 1.710 11.310 2.505 ;
        RECT  10.780 1.080 11.120 1.420 ;
        RECT  10.970 1.710 11.080 2.050 ;
        RECT  9.785 1.765 10.970 1.995 ;
        RECT  10.620 2.955 10.960 3.440 ;
        RECT  10.305 2.225 10.640 2.455 ;
        RECT  10.075 2.225 10.305 3.785 ;
        RECT  8.860 3.555 10.075 3.785 ;
        RECT  9.555 1.765 9.785 3.265 ;
        RECT  9.040 1.765 9.555 1.995 ;
        RECT  9.060 3.035 9.555 3.265 ;
        RECT  8.970 2.270 9.310 2.610 ;
        RECT  8.720 2.980 9.060 3.320 ;
        RECT  8.885 1.160 9.040 1.995 ;
        RECT  8.375 2.325 8.970 2.555 ;
        RECT  8.755 0.630 8.885 1.995 ;
        RECT  8.520 3.555 8.860 4.010 ;
        RECT  8.655 0.630 8.755 1.500 ;
        RECT  8.605 0.630 8.655 0.970 ;
        RECT  6.205 3.555 8.520 3.785 ;
        RECT  8.200 1.145 8.375 3.210 ;
        RECT  8.145 0.960 8.200 3.210 ;
        RECT  7.860 0.960 8.145 1.375 ;
        RECT  7.740 2.980 8.145 3.210 ;
        RECT  7.490 1.605 7.830 1.945 ;
        RECT  7.400 2.980 7.740 3.320 ;
        RECT  5.750 1.605 7.490 1.835 ;
        RECT  6.965 2.980 7.400 3.210 ;
        RECT  6.735 2.175 6.965 3.210 ;
        RECT  6.640 2.175 6.735 2.405 ;
        RECT  6.300 2.065 6.640 2.405 ;
        RECT  5.975 3.555 6.205 4.285 ;
        RECT  5.285 4.055 5.975 4.285 ;
        RECT  5.745 1.095 5.750 1.835 ;
        RECT  5.560 1.095 5.745 3.720 ;
        RECT  5.515 1.040 5.560 3.720 ;
        RECT  5.220 1.040 5.515 1.380 ;
        RECT  5.280 1.665 5.285 4.285 ;
        RECT  5.055 1.610 5.280 4.285 ;
        RECT  4.940 1.610 5.055 1.950 ;
        RECT  4.360 2.910 5.055 3.140 ;
        RECT  4.595 3.380 4.825 3.910 ;
        RECT  4.420 0.775 4.760 1.115 ;
        RECT  2.980 3.680 4.595 3.910 ;
        RECT  2.660 0.860 4.420 1.090 ;
        RECT  4.130 2.910 4.360 3.450 ;
        RECT  2.520 3.220 4.130 3.450 ;
        RECT  2.415 1.360 3.680 1.590 ;
        RECT  2.750 3.680 2.980 4.025 ;
        RECT  1.850 3.795 2.750 4.025 ;
        RECT  2.430 0.650 2.660 1.090 ;
        RECT  2.290 3.220 2.520 3.565 ;
        RECT  2.415 2.650 2.470 2.990 ;
        RECT  1.700 0.650 2.430 0.880 ;
        RECT  2.185 1.360 2.415 2.990 ;
        RECT  0.600 3.335 2.290 3.565 ;
        RECT  1.640 1.360 2.185 1.590 ;
        RECT  2.130 2.650 2.185 2.990 ;
        RECT  1.940 2.760 2.130 2.990 ;
        RECT  1.600 2.760 1.940 3.105 ;
        RECT  0.380 1.255 0.600 1.595 ;
        RECT  0.380 2.960 0.600 3.565 ;
        RECT  0.370 1.255 0.380 3.565 ;
        RECT  0.150 1.255 0.370 3.300 ;
    END
END SDFFSX4

MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.990 3.995 12.400 4.340 ;
        RECT  11.130 3.995 11.990 4.225 ;
        RECT  10.900 3.995 11.130 4.310 ;
        RECT  10.080 4.080 10.900 4.310 ;
        RECT  9.850 4.005 10.080 4.310 ;
        RECT  7.140 4.005 9.850 4.235 ;
        RECT  6.910 4.005 7.140 4.240 ;
        RECT  6.855 4.010 6.910 4.240 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.995 3.305 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.820 1.655 2.100 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.830 1.240 14.965 1.515 ;
        RECT  14.600 0.685 14.830 2.970 ;
        RECT  14.290 0.685 14.600 0.915 ;
        RECT  14.500 2.740 14.600 2.970 ;
        RECT  14.160 2.740 14.500 3.080 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.070 1.325 16.285 3.145 ;
        RECT  16.055 0.745 16.070 3.145 ;
        RECT  15.730 0.745 16.055 1.555 ;
        RECT  15.940 2.915 16.055 3.220 ;
        RECT  15.600 2.915 15.940 4.195 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.170 1.820 4.510 2.500 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.830 0.820 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.295 -0.400 16.500 0.400 ;
        RECT  15.065 -0.400 15.295 1.005 ;
        RECT  13.370 -0.400 15.065 0.400 ;
        RECT  13.030 -0.400 13.370 0.575 ;
        RECT  11.550 -0.400 13.030 0.400 ;
        RECT  11.210 -0.400 11.550 1.095 ;
        RECT  9.005 -0.400 11.210 0.400 ;
        RECT  8.775 -0.400 9.005 1.440 ;
        RECT  6.780 -0.400 8.775 0.400 ;
        RECT  6.440 -0.400 6.780 1.130 ;
        RECT  3.585 -0.400 6.440 0.400 ;
        RECT  3.245 -0.400 3.585 0.575 ;
        RECT  1.425 -0.400 3.245 0.400 ;
        RECT  1.085 -0.400 1.425 0.575 ;
        RECT  0.000 -0.400 1.085 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.220 4.640 16.500 5.440 ;
        RECT  14.880 3.895 15.220 5.440 ;
        RECT  13.240 4.640 14.880 5.440 ;
        RECT  12.900 3.445 13.240 5.440 ;
        RECT  11.760 4.640 12.900 5.440 ;
        RECT  11.420 4.465 11.760 5.440 ;
        RECT  9.495 4.640 11.420 5.440 ;
        RECT  8.940 4.465 9.495 5.440 ;
        RECT  8.020 4.640 8.940 5.440 ;
        RECT  7.680 4.465 8.020 5.440 ;
        RECT  6.620 4.640 7.680 5.440 ;
        RECT  6.280 4.465 6.620 5.440 ;
        RECT  3.540 4.640 6.280 5.440 ;
        RECT  3.200 3.955 3.540 5.440 ;
        RECT  1.080 4.640 3.200 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.370 2.070 15.590 2.410 ;
        RECT  15.140 2.070 15.370 3.545 ;
        RECT  13.960 3.315 15.140 3.545 ;
        RECT  13.930 1.345 14.090 1.685 ;
        RECT  13.930 3.315 13.960 3.785 ;
        RECT  13.700 1.345 13.930 3.785 ;
        RECT  13.620 3.445 13.700 3.785 ;
        RECT  13.325 2.015 13.435 2.355 ;
        RECT  13.095 1.325 13.325 3.170 ;
        RECT  12.830 1.325 13.095 1.555 ;
        RECT  12.520 2.940 13.095 3.170 ;
        RECT  12.490 1.260 12.830 1.600 ;
        RECT  12.655 2.190 12.760 2.530 ;
        RECT  12.420 2.190 12.655 2.670 ;
        RECT  12.180 2.940 12.520 3.750 ;
        RECT  11.245 1.325 12.490 1.555 ;
        RECT  10.545 2.440 12.420 2.670 ;
        RECT  11.015 1.325 11.245 2.205 ;
        RECT  10.905 1.865 11.015 2.205 ;
        RECT  10.545 1.360 10.550 1.700 ;
        RECT  10.315 1.360 10.545 3.850 ;
        RECT  10.210 1.360 10.315 1.700 ;
        RECT  9.835 2.540 10.065 3.775 ;
        RECT  9.550 1.870 9.980 2.210 ;
        RECT  6.245 3.545 9.835 3.775 ;
        RECT  9.320 1.670 9.550 3.020 ;
        RECT  8.545 1.670 9.320 1.900 ;
        RECT  8.780 2.790 9.320 3.020 ;
        RECT  8.085 2.140 9.090 2.480 ;
        RECT  8.440 2.790 8.780 3.130 ;
        RECT  8.315 0.725 8.545 1.900 ;
        RECT  7.530 0.725 8.315 0.955 ;
        RECT  7.855 1.440 8.085 3.230 ;
        RECT  6.460 3.000 7.855 3.230 ;
        RECT  6.930 2.445 7.570 2.675 ;
        RECT  7.190 0.635 7.530 0.955 ;
        RECT  6.700 1.945 6.930 2.675 ;
        RECT  5.690 1.945 6.700 2.175 ;
        RECT  6.230 2.415 6.460 3.230 ;
        RECT  6.015 3.545 6.245 4.085 ;
        RECT  6.120 2.415 6.230 2.755 ;
        RECT  5.475 3.855 6.015 4.085 ;
        RECT  5.690 0.760 5.745 1.100 ;
        RECT  5.460 0.760 5.690 3.285 ;
        RECT  5.245 3.855 5.475 4.405 ;
        RECT  5.405 0.760 5.460 1.100 ;
        RECT  5.215 2.945 5.460 3.285 ;
        RECT  4.985 4.175 5.245 4.405 ;
        RECT  4.985 1.505 5.170 1.955 ;
        RECT  4.755 1.505 4.985 4.405 ;
        RECT  4.605 0.760 4.945 1.100 ;
        RECT  4.000 4.175 4.755 4.405 ;
        RECT  2.640 0.815 4.605 1.045 ;
        RECT  4.245 3.035 4.475 3.945 ;
        RECT  2.425 3.035 4.245 3.265 ;
        RECT  3.770 3.495 4.000 4.405 ;
        RECT  3.525 1.295 3.865 1.635 ;
        RECT  2.970 3.495 3.770 3.725 ;
        RECT  2.470 1.350 3.525 1.580 ;
        RECT  2.740 3.495 2.970 4.365 ;
        RECT  1.685 4.135 2.740 4.365 ;
        RECT  2.410 0.695 2.640 1.045 ;
        RECT  2.240 1.350 2.470 2.755 ;
        RECT  2.195 3.035 2.425 3.900 ;
        RECT  1.885 0.695 2.410 0.925 ;
        RECT  1.885 1.350 2.240 1.690 ;
        RECT  2.130 2.415 2.240 2.755 ;
        RECT  2.040 3.560 2.195 3.900 ;
        RECT  1.880 2.525 2.130 2.755 ;
        RECT  1.650 2.525 1.880 3.160 ;
        RECT  1.455 3.595 1.685 4.365 ;
        RECT  1.540 2.820 1.650 3.160 ;
        RECT  1.280 3.595 1.455 3.825 ;
        RECT  1.050 2.350 1.280 3.825 ;
        RECT  0.410 2.350 1.050 2.580 ;
        RECT  0.520 3.540 1.050 3.825 ;
        RECT  0.410 1.230 0.520 1.570 ;
        RECT  0.180 3.485 0.520 3.825 ;
        RECT  0.180 1.230 0.410 2.580 ;
    END
END SDFFSX2

MACRO SDFFSX1
    CLASS CORE ;
    FOREIGN SDFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.020 4.060 12.650 4.410 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.750 2.110 3.335 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.830 1.815 1.600 2.100 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.200 0.865 14.430 3.950 ;
        RECT  13.620 0.865 14.200 1.095 ;
        RECT  13.960 3.720 14.200 3.950 ;
        RECT  13.645 3.720 13.960 4.105 ;
        RECT  13.415 3.720 13.645 4.315 ;
        RECT  13.280 0.700 13.620 1.095 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.200 2.855 15.540 3.665 ;
        RECT  15.040 1.250 15.380 1.590 ;
        RECT  15.040 2.855 15.200 3.220 ;
        RECT  14.965 1.285 15.040 1.590 ;
        RECT  14.965 2.635 15.040 3.220 ;
        RECT  14.735 1.360 14.965 3.085 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.510 2.375 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.830 0.755 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.570 -0.400 15.840 0.400 ;
        RECT  14.230 -0.400 14.570 0.575 ;
        RECT  12.800 -0.400 14.230 0.400 ;
        RECT  12.460 -0.400 12.800 0.575 ;
        RECT  11.400 -0.400 12.460 0.400 ;
        RECT  11.060 -0.400 11.400 0.575 ;
        RECT  9.005 -0.400 11.060 0.400 ;
        RECT  8.775 -0.400 9.005 1.010 ;
        RECT  6.980 -0.400 8.775 0.400 ;
        RECT  6.640 -0.400 6.980 1.050 ;
        RECT  3.585 -0.400 6.640 0.400 ;
        RECT  3.245 -0.400 3.585 0.575 ;
        RECT  1.425 -0.400 3.245 0.400 ;
        RECT  1.085 -0.400 1.425 0.575 ;
        RECT  0.000 -0.400 1.085 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.705 4.640 15.840 5.440 ;
        RECT  14.305 4.465 14.705 5.440 ;
        RECT  13.110 4.640 14.305 5.440 ;
        RECT  13.110 2.920 13.240 3.260 ;
        RECT  12.880 2.920 13.110 5.440 ;
        RECT  11.790 4.640 12.880 5.440 ;
        RECT  11.450 4.140 11.790 5.440 ;
        RECT  9.280 4.640 11.450 5.440 ;
        RECT  8.940 4.140 9.280 5.440 ;
        RECT  8.020 4.640 8.940 5.440 ;
        RECT  7.680 4.140 8.020 5.440 ;
        RECT  6.620 4.640 7.680 5.440 ;
        RECT  6.280 4.465 6.620 5.440 ;
        RECT  3.485 4.640 6.280 5.440 ;
        RECT  3.255 4.100 3.485 5.440 ;
        RECT  1.080 4.640 3.255 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.905 1.550 13.970 2.745 ;
        RECT  13.740 1.550 13.905 3.260 ;
        RECT  13.660 1.550 13.740 1.780 ;
        RECT  13.675 2.515 13.740 3.260 ;
        RECT  13.320 1.440 13.660 1.780 ;
        RECT  12.520 2.025 13.355 2.255 ;
        RECT  12.290 1.540 12.520 3.400 ;
        RECT  11.740 1.540 12.290 1.770 ;
        RECT  12.180 3.060 12.290 3.400 ;
        RECT  11.700 2.380 12.040 2.720 ;
        RECT  11.400 1.430 11.740 1.770 ;
        RECT  10.545 2.435 11.700 2.665 ;
        RECT  11.050 1.430 11.400 1.660 ;
        RECT  10.815 1.160 11.050 1.660 ;
        RECT  10.710 1.160 10.815 1.500 ;
        RECT  10.545 3.410 10.600 3.750 ;
        RECT  10.325 1.875 10.545 3.750 ;
        RECT  10.315 1.435 10.325 3.750 ;
        RECT  10.095 1.435 10.315 2.105 ;
        RECT  10.260 3.410 10.315 3.750 ;
        RECT  9.890 4.020 10.230 4.360 ;
        RECT  9.965 1.435 10.095 1.780 ;
        RECT  9.910 1.440 9.965 1.780 ;
        RECT  9.775 2.335 9.940 2.675 ;
        RECT  9.740 4.020 9.890 4.250 ;
        RECT  9.680 2.335 9.775 3.145 ;
        RECT  9.510 3.670 9.740 4.250 ;
        RECT  9.450 1.245 9.680 3.145 ;
        RECT  6.245 3.670 9.510 3.900 ;
        RECT  8.545 1.245 9.450 1.475 ;
        RECT  8.725 2.915 9.450 3.145 ;
        RECT  8.875 2.165 9.215 2.505 ;
        RECT  8.265 2.220 8.875 2.450 ;
        RECT  8.495 2.915 8.725 3.420 ;
        RECT  8.315 0.725 8.545 1.475 ;
        RECT  8.035 0.725 8.315 0.955 ;
        RECT  8.085 2.220 8.265 3.310 ;
        RECT  8.035 1.420 8.085 3.310 ;
        RECT  7.805 0.675 8.035 0.955 ;
        RECT  7.855 1.420 8.035 2.450 ;
        RECT  7.420 3.080 8.035 3.310 ;
        RECT  7.310 0.675 7.805 0.905 ;
        RECT  7.460 2.445 7.570 2.785 ;
        RECT  7.230 2.180 7.460 2.785 ;
        RECT  7.080 3.080 7.420 3.420 ;
        RECT  5.690 2.180 7.230 2.410 ;
        RECT  6.460 3.080 7.080 3.310 ;
        RECT  6.230 2.640 6.460 3.310 ;
        RECT  6.015 3.670 6.245 4.085 ;
        RECT  6.120 2.640 6.230 2.980 ;
        RECT  5.685 3.855 6.015 4.085 ;
        RECT  5.690 0.760 5.745 1.100 ;
        RECT  5.460 0.760 5.690 3.125 ;
        RECT  5.400 3.855 5.685 4.405 ;
        RECT  5.405 0.760 5.460 1.100 ;
        RECT  5.445 2.895 5.460 3.125 ;
        RECT  5.215 2.895 5.445 3.520 ;
        RECT  4.985 4.175 5.400 4.405 ;
        RECT  5.000 1.400 5.230 2.430 ;
        RECT  4.985 2.200 5.000 2.430 ;
        RECT  4.755 2.200 4.985 4.405 ;
        RECT  4.655 0.815 4.945 1.045 ;
        RECT  3.945 4.175 4.755 4.405 ;
        RECT  4.425 0.815 4.655 1.095 ;
        RECT  4.415 3.605 4.525 3.945 ;
        RECT  2.640 0.865 4.425 1.095 ;
        RECT  4.185 3.035 4.415 3.945 ;
        RECT  2.380 3.035 4.185 3.265 ;
        RECT  3.715 3.630 3.945 4.405 ;
        RECT  3.525 1.350 3.865 1.690 ;
        RECT  3.020 3.630 3.715 3.860 ;
        RECT  2.415 1.460 3.525 1.690 ;
        RECT  2.790 3.630 3.020 4.365 ;
        RECT  1.685 4.135 2.790 4.365 ;
        RECT  2.410 0.695 2.640 1.095 ;
        RECT  2.415 2.465 2.470 2.805 ;
        RECT  2.225 1.460 2.415 2.805 ;
        RECT  1.885 0.695 2.410 0.925 ;
        RECT  2.150 3.035 2.380 3.900 ;
        RECT  2.185 1.350 2.225 2.805 ;
        RECT  1.885 1.350 2.185 1.690 ;
        RECT  2.130 2.465 2.185 2.805 ;
        RECT  2.040 3.560 2.150 3.900 ;
        RECT  1.880 2.575 2.130 2.805 ;
        RECT  1.650 2.575 1.880 3.160 ;
        RECT  1.455 3.650 1.685 4.365 ;
        RECT  1.540 2.820 1.650 3.160 ;
        RECT  1.215 3.650 1.455 3.880 ;
        RECT  0.985 2.350 1.215 3.880 ;
        RECT  0.410 2.350 0.985 2.580 ;
        RECT  0.180 3.540 0.985 3.880 ;
        RECT  0.410 1.190 0.520 1.530 ;
        RECT  0.180 1.190 0.410 2.580 ;
    END
END SDFFSX1

MACRO SDFFRHQXL
    CLASS CORE ;
    FOREIGN SDFFRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.290 2.380 3.745 2.635 ;
        RECT  3.005 2.050 3.290 2.635 ;
        RECT  2.950 2.050 3.005 2.390 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 1.820 1.870 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.950 2.965 14.965 3.195 ;
        RECT  14.160 2.910 14.950 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.360 1.270 16.375 3.195 ;
        RECT  16.145 1.270 16.360 4.055 ;
        RECT  15.290 1.270 16.145 1.500 ;
        RECT  16.055 2.965 16.145 4.055 ;
        RECT  15.960 3.715 16.055 4.055 ;
        RECT  15.060 0.700 15.290 1.500 ;
        RECT  14.950 0.700 15.060 1.040 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 1.750 4.480 2.110 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.170 1.105 2.635 ;
        RECT  0.630 2.170 0.875 2.625 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.090 -0.400 16.500 0.400 ;
        RECT  15.750 -0.400 16.090 1.040 ;
        RECT  14.485 -0.400 15.750 0.400 ;
        RECT  13.545 -0.400 14.485 0.575 ;
        RECT  12.405 -0.400 13.545 0.400 ;
        RECT  12.065 -0.400 12.405 0.575 ;
        RECT  9.430 -0.400 12.065 0.400 ;
        RECT  9.090 -0.400 9.430 1.160 ;
        RECT  6.740 -0.400 9.090 0.400 ;
        RECT  8.040 1.460 8.150 1.800 ;
        RECT  7.810 1.145 8.040 1.800 ;
        RECT  6.740 1.145 7.810 1.375 ;
        RECT  6.400 -0.400 6.740 1.375 ;
        RECT  3.255 -0.400 6.400 0.400 ;
        RECT  2.915 -0.400 3.255 0.575 ;
        RECT  1.130 -0.400 2.915 0.400 ;
        RECT  0.790 -0.400 1.130 0.575 ;
        RECT  0.000 -0.400 0.790 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.020 4.640 16.500 5.440 ;
        RECT  14.680 3.505 15.020 5.440 ;
        RECT  13.920 3.505 14.680 3.735 ;
        RECT  12.730 4.640 14.680 5.440 ;
        RECT  13.690 3.140 13.920 3.735 ;
        RECT  13.580 3.140 13.690 3.480 ;
        RECT  12.315 4.465 12.730 5.440 ;
        RECT  9.770 4.640 12.315 5.440 ;
        RECT  9.430 4.465 9.770 5.440 ;
        RECT  6.680 4.640 9.430 5.440 ;
        RECT  6.340 4.000 6.680 5.440 ;
        RECT  3.500 4.640 6.340 5.440 ;
        RECT  3.160 4.130 3.500 5.440 ;
        RECT  0.920 4.640 3.160 5.440 ;
        RECT  0.580 3.835 0.920 5.440 ;
        RECT  0.000 4.640 0.580 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.440 1.765 15.820 1.995 ;
        RECT  13.805 2.440 15.255 2.670 ;
        RECT  14.210 0.865 14.440 1.995 ;
        RECT  13.265 3.965 14.220 4.195 ;
        RECT  12.765 0.865 14.210 1.095 ;
        RECT  13.805 1.375 13.885 1.715 ;
        RECT  13.775 1.375 13.805 2.670 ;
        RECT  13.545 1.375 13.775 2.680 ;
        RECT  13.265 2.210 13.545 2.680 ;
        RECT  13.225 2.210 13.265 4.195 ;
        RECT  13.035 2.405 13.225 4.195 ;
        RECT  12.745 1.410 13.085 1.750 ;
        RECT  8.425 3.965 13.035 4.195 ;
        RECT  12.395 0.865 12.765 1.145 ;
        RECT  12.680 1.520 12.745 1.750 ;
        RECT  12.450 1.520 12.680 3.445 ;
        RECT  12.260 2.540 12.450 3.445 ;
        RECT  11.865 0.865 12.395 1.095 ;
        RECT  12.095 2.540 12.260 2.890 ;
        RECT  11.635 0.865 11.865 3.600 ;
        RECT  11.040 0.865 11.635 1.105 ;
        RECT  11.310 3.370 11.635 3.600 ;
        RECT  11.120 1.610 11.320 1.950 ;
        RECT  10.970 3.370 11.310 3.710 ;
        RECT  10.890 1.610 11.120 3.055 ;
        RECT  10.700 0.865 11.040 1.285 ;
        RECT  10.590 1.595 10.660 3.655 ;
        RECT  10.455 1.595 10.590 3.710 ;
        RECT  10.430 1.045 10.455 3.710 ;
        RECT  10.240 1.045 10.430 1.825 ;
        RECT  10.250 3.370 10.430 3.710 ;
        RECT  10.225 0.990 10.240 1.825 ;
        RECT  9.900 0.990 10.225 1.330 ;
        RECT  9.975 2.280 10.200 2.620 ;
        RECT  9.745 1.630 9.975 3.480 ;
        RECT  9.010 1.630 9.745 1.860 ;
        RECT  9.270 3.250 9.745 3.480 ;
        RECT  9.405 2.575 9.515 2.915 ;
        RECT  9.175 2.205 9.405 2.915 ;
        RECT  8.930 3.250 9.270 3.590 ;
        RECT  7.505 2.205 9.175 2.435 ;
        RECT  8.845 1.520 9.010 1.860 ;
        RECT  8.615 0.685 8.845 1.860 ;
        RECT  7.000 0.685 8.615 0.915 ;
        RECT  8.195 2.680 8.425 4.195 ;
        RECT  7.960 2.680 8.195 3.020 ;
        RECT  7.275 1.635 7.505 3.680 ;
        RECT  6.335 1.635 7.275 1.895 ;
        RECT  7.050 3.340 7.275 3.680 ;
        RECT  6.705 2.635 7.045 2.985 ;
        RECT  5.575 2.755 6.705 2.985 ;
        RECT  6.105 1.635 6.335 2.370 ;
        RECT  5.995 2.030 6.105 2.370 ;
        RECT  5.470 3.740 5.810 4.080 ;
        RECT  5.435 0.950 5.575 2.985 ;
        RECT  4.945 3.740 5.470 3.970 ;
        RECT  5.345 0.950 5.435 3.325 ;
        RECT  5.340 0.950 5.345 1.180 ;
        RECT  5.205 2.715 5.345 3.325 ;
        RECT  5.000 0.840 5.340 1.180 ;
        RECT  4.715 1.655 4.945 3.970 ;
        RECT  2.360 3.075 4.715 3.305 ;
        RECT  4.280 0.820 4.620 1.160 ;
        RECT  4.255 3.595 4.485 4.185 ;
        RECT  1.905 0.875 4.280 1.105 ;
        RECT  2.835 3.595 4.255 3.825 ;
        RECT  3.200 1.375 3.540 1.715 ;
        RECT  2.360 1.485 3.200 1.715 ;
        RECT  2.605 3.595 2.835 4.060 ;
        RECT  2.000 3.830 2.605 4.060 ;
        RECT  2.360 2.500 2.590 2.840 ;
        RECT  2.130 1.460 2.360 2.840 ;
        RECT  2.130 3.075 2.360 3.600 ;
        RECT  1.840 2.610 2.130 2.840 ;
        RECT  1.215 3.370 2.130 3.600 ;
        RECT  1.675 0.630 1.905 1.105 ;
        RECT  1.610 2.610 1.840 3.140 ;
        RECT  1.490 0.630 1.675 0.860 ;
        RECT  1.500 2.800 1.610 3.140 ;
        RECT  0.985 2.890 1.215 3.600 ;
        RECT  0.520 2.890 0.985 3.120 ;
        RECT  0.395 1.400 0.520 1.740 ;
        RECT  0.395 2.855 0.520 3.120 ;
        RECT  0.165 1.400 0.395 3.120 ;
    END
END SDFFRHQXL

MACRO SDFFRHQX4
    CLASS CORE ;
    FOREIGN SDFFRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRHQXL ;
    SIZE 24.420 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.820 3.160 3.385 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 2.360 4.160 2.590 ;
        RECT  3.515 2.360 3.745 2.635 ;
        RECT  3.165 2.360 3.515 2.590 ;
        RECT  2.935 1.905 3.165 2.590 ;
        RECT  2.630 1.905 2.935 2.135 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.280 1.835 18.265 2.100 ;
        RECT  17.275 1.835 17.280 2.065 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.110 2.970 24.165 3.910 ;
        RECT  23.825 2.965 24.110 3.910 ;
        RECT  23.620 2.965 23.825 3.220 ;
        RECT  23.240 1.465 23.620 3.220 ;
        RECT  22.920 1.465 23.240 1.695 ;
        RECT  21.605 2.990 23.240 3.220 ;
        RECT  22.580 0.750 22.920 1.695 ;
        RECT  21.480 1.465 22.580 1.695 ;
        RECT  21.265 2.970 21.605 3.910 ;
        RECT  21.195 0.750 21.480 1.695 ;
        RECT  21.140 0.750 21.195 1.690 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 2.965 4.600 3.325 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.000 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.640 -0.400 24.420 0.400 ;
        RECT  23.300 -0.400 23.640 1.050 ;
        RECT  22.200 -0.400 23.300 0.400 ;
        RECT  21.860 -0.400 22.200 1.050 ;
        RECT  20.515 -0.400 21.860 0.400 ;
        RECT  20.285 -0.400 20.515 1.575 ;
        RECT  18.785 -0.400 20.285 0.400 ;
        RECT  18.445 -0.400 18.785 0.575 ;
        RECT  17.305 -0.400 18.445 0.400 ;
        RECT  16.965 -0.400 17.305 1.190 ;
        RECT  11.765 -0.400 16.965 0.400 ;
        RECT  11.425 -0.400 11.765 1.320 ;
        RECT  10.325 -0.400 11.425 0.400 ;
        RECT  9.985 -0.400 10.325 1.490 ;
        RECT  8.650 -0.400 9.985 0.400 ;
        RECT  8.650 1.260 8.705 1.600 ;
        RECT  8.420 -0.400 8.650 1.600 ;
        RECT  7.225 -0.400 8.420 0.400 ;
        RECT  8.365 1.260 8.420 1.600 ;
        RECT  6.885 -0.400 7.225 0.970 ;
        RECT  4.010 -0.400 6.885 0.400 ;
        RECT  3.670 -0.400 4.010 0.575 ;
        RECT  1.285 -0.400 3.670 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.885 4.640 24.420 5.440 ;
        RECT  22.545 3.760 22.885 5.440 ;
        RECT  20.270 4.640 22.545 5.440 ;
        RECT  20.040 3.055 20.270 5.440 ;
        RECT  18.625 4.640 20.040 5.440 ;
        RECT  18.285 4.465 18.625 5.440 ;
        RECT  16.980 4.640 18.285 5.440 ;
        RECT  16.640 4.090 16.980 5.440 ;
        RECT  11.985 4.640 16.640 5.440 ;
        RECT  11.645 4.465 11.985 5.440 ;
        RECT  10.460 4.640 11.645 5.440 ;
        RECT  10.230 4.060 10.460 5.440 ;
        RECT  9.035 4.640 10.230 5.440 ;
        RECT  8.695 4.465 9.035 5.440 ;
        RECT  7.145 4.640 8.695 5.440 ;
        RECT  6.805 4.465 7.145 5.440 ;
        RECT  1.320 4.640 6.805 5.440 ;
        RECT  0.980 4.465 1.320 5.440 ;
        RECT  0.000 4.640 0.980 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.275 2.125 22.520 2.355 ;
        RECT  20.055 2.125 20.275 2.495 ;
        RECT  19.825 0.805 20.055 2.495 ;
        RECT  18.025 0.805 19.825 1.035 ;
        RECT  19.810 2.265 19.825 2.495 ;
        RECT  19.580 2.265 19.810 4.175 ;
        RECT  19.365 1.265 19.595 1.775 ;
        RECT  17.450 3.945 19.580 4.175 ;
        RECT  18.865 1.545 19.365 1.775 ;
        RECT  19.120 2.200 19.350 3.715 ;
        RECT  17.960 3.485 19.120 3.715 ;
        RECT  18.635 1.545 18.865 3.255 ;
        RECT  17.045 2.565 18.635 2.795 ;
        RECT  17.740 0.805 18.025 1.330 ;
        RECT  17.730 3.155 17.960 3.715 ;
        RECT  17.685 0.990 17.740 1.330 ;
        RECT  16.580 3.155 17.730 3.385 ;
        RECT  17.220 3.620 17.450 4.175 ;
        RECT  16.375 3.620 17.220 3.850 ;
        RECT  16.815 2.200 17.045 2.795 ;
        RECT  16.225 2.200 16.815 2.430 ;
        RECT  16.350 2.725 16.580 3.385 ;
        RECT  16.145 3.620 16.375 4.365 ;
        RECT  15.810 2.725 16.350 2.955 ;
        RECT  12.445 4.135 16.145 4.365 ;
        RECT  15.810 1.100 15.945 1.440 ;
        RECT  15.685 3.200 15.915 3.845 ;
        RECT  15.580 0.675 15.810 2.955 ;
        RECT  13.025 3.615 15.685 3.845 ;
        RECT  14.505 0.675 15.580 0.905 ;
        RECT  15.300 2.635 15.580 2.955 ;
        RECT  14.065 2.635 15.300 2.865 ;
        RECT  14.970 1.195 15.225 1.425 ;
        RECT  14.740 1.195 14.970 1.925 ;
        RECT  13.540 3.095 14.880 3.325 ;
        RECT  13.785 1.695 14.740 1.925 ;
        RECT  14.165 0.675 14.505 1.380 ;
        RECT  12.685 0.675 14.165 0.905 ;
        RECT  13.835 2.520 14.065 2.865 ;
        RECT  13.540 1.195 13.785 1.925 ;
        RECT  13.310 1.195 13.540 3.325 ;
        RECT  13.235 1.195 13.310 1.925 ;
        RECT  13.255 2.905 13.310 3.325 ;
        RECT  11.895 2.905 13.255 3.135 ;
        RECT  12.430 1.195 13.235 1.425 ;
        RECT  12.795 3.425 13.025 3.845 ;
        RECT  12.730 1.770 12.960 2.435 ;
        RECT  11.380 3.425 12.795 3.655 ;
        RECT  11.380 2.205 12.730 2.435 ;
        RECT  12.215 4.005 12.445 4.365 ;
        RECT  12.200 1.195 12.430 1.785 ;
        RECT  10.920 4.005 12.215 4.235 ;
        RECT  11.045 1.555 12.200 1.785 ;
        RECT  11.665 2.770 11.895 3.135 ;
        RECT  11.150 2.205 11.380 3.655 ;
        RECT  10.395 2.205 11.150 2.435 ;
        RECT  10.815 1.135 11.045 1.785 ;
        RECT  10.690 3.395 10.920 4.235 ;
        RECT  10.705 1.135 10.815 1.475 ;
        RECT  9.785 3.395 10.690 3.625 ;
        RECT  10.395 2.750 10.450 3.090 ;
        RECT  10.165 1.775 10.395 3.090 ;
        RECT  9.600 1.775 10.165 2.005 ;
        RECT  10.110 2.750 10.165 3.090 ;
        RECT  9.700 3.860 9.930 4.220 ;
        RECT  9.555 2.295 9.785 3.625 ;
        RECT  8.805 3.860 9.700 4.090 ;
        RECT  9.490 1.260 9.600 2.005 ;
        RECT  8.305 2.295 9.555 2.525 ;
        RECT  9.370 0.675 9.490 2.005 ;
        RECT  9.260 0.675 9.370 1.600 ;
        RECT  8.075 2.935 9.320 3.325 ;
        RECT  8.895 0.675 9.260 0.905 ;
        RECT  8.575 3.860 8.805 4.175 ;
        RECT  6.195 3.945 8.575 4.175 ;
        RECT  7.845 1.235 8.075 3.325 ;
        RECT  7.700 1.235 7.845 1.600 ;
        RECT  7.835 2.930 7.845 3.325 ;
        RECT  7.340 2.930 7.835 3.270 ;
        RECT  7.250 2.015 7.605 2.585 ;
        RECT  6.925 2.930 7.340 3.160 ;
        RECT  6.165 2.015 7.250 2.245 ;
        RECT  6.695 2.570 6.925 3.160 ;
        RECT  6.585 2.570 6.695 2.910 ;
        RECT  6.195 2.730 6.250 3.070 ;
        RECT  5.965 2.730 6.195 4.175 ;
        RECT  6.000 2.015 6.165 2.365 ;
        RECT  6.000 0.900 6.055 1.240 ;
        RECT  5.770 0.900 6.000 2.365 ;
        RECT  5.910 2.730 5.965 3.070 ;
        RECT  5.060 3.670 5.965 3.915 ;
        RECT  5.715 0.900 5.770 1.240 ;
        RECT  5.665 2.135 5.770 2.365 ;
        RECT  5.435 2.135 5.665 3.435 ;
        RECT  5.290 1.470 5.520 1.835 ;
        RECT  4.995 0.875 5.345 1.155 ;
        RECT  5.060 1.605 5.290 1.835 ;
        RECT  4.830 1.605 5.060 3.915 ;
        RECT  2.650 0.875 4.995 1.105 ;
        RECT  2.080 4.145 4.960 4.375 ;
        RECT  2.545 3.685 4.830 3.915 ;
        RECT  3.820 1.445 4.160 1.810 ;
        RECT  2.020 1.445 3.820 1.675 ;
        RECT  2.310 0.875 2.650 1.205 ;
        RECT  2.315 3.255 2.545 3.915 ;
        RECT  0.520 3.255 2.315 3.485 ;
        RECT  1.850 3.715 2.080 4.375 ;
        RECT  2.020 2.000 2.075 2.340 ;
        RECT  1.790 1.075 2.020 3.025 ;
        RECT  1.720 3.715 1.850 3.945 ;
        RECT  1.610 1.075 1.790 1.305 ;
        RECT  1.735 2.000 1.790 2.340 ;
        RECT  1.680 2.795 1.790 3.025 ;
        RECT  0.395 0.700 0.520 1.510 ;
        RECT  0.395 3.060 0.520 4.000 ;
        RECT  0.165 0.700 0.395 4.000 ;
    END
END SDFFRHQX4

MACRO SDFFRHQX2
    CLASS CORE ;
    FOREIGN SDFFRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRHQXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.295 2.380 3.745 2.640 ;
        RECT  2.955 2.300 3.295 2.640 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.745 1.870 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.055 2.655 16.590 3.205 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.800 1.155 19.030 3.060 ;
        RECT  17.680 1.155 18.800 1.385 ;
        RECT  18.340 2.830 18.800 3.060 ;
        RECT  18.000 2.830 18.340 4.030 ;
        RECT  17.670 0.945 17.680 1.385 ;
        RECT  17.330 0.635 17.670 1.445 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 1.755 4.480 2.140 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.125 1.180 2.590 ;
        RECT  0.875 2.125 1.105 2.635 ;
        RECT  0.600 2.125 0.875 2.590 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.430 -0.400 19.800 0.400 ;
        RECT  18.090 -0.400 18.430 0.575 ;
        RECT  16.685 -0.400 18.090 0.400 ;
        RECT  15.745 -0.400 16.685 0.575 ;
        RECT  14.400 -0.400 15.745 0.400 ;
        RECT  14.060 -0.400 14.400 0.575 ;
        RECT  10.485 -0.400 14.060 0.400 ;
        RECT  10.145 -0.400 10.485 1.290 ;
        RECT  6.590 -0.400 10.145 0.400 ;
        RECT  7.750 1.210 8.090 1.570 ;
        RECT  6.590 1.210 7.750 1.440 ;
        RECT  6.360 -0.400 6.590 1.440 ;
        RECT  6.250 -0.400 6.360 1.435 ;
        RECT  3.145 -0.400 6.250 0.400 ;
        RECT  2.805 -0.400 3.145 0.575 ;
        RECT  1.080 -0.400 2.805 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 4.640 19.800 5.440 ;
        RECT  19.280 3.295 19.620 5.440 ;
        RECT  16.970 4.640 19.280 5.440 ;
        RECT  16.630 4.465 16.970 5.440 ;
        RECT  15.570 4.640 16.630 5.440 ;
        RECT  15.230 4.465 15.570 5.440 ;
        RECT  14.385 4.640 15.230 5.440 ;
        RECT  13.945 4.465 14.385 5.440 ;
        RECT  10.505 4.640 13.945 5.440 ;
        RECT  10.165 4.465 10.505 5.440 ;
        RECT  6.680 4.640 10.165 5.440 ;
        RECT  6.340 4.125 6.680 5.440 ;
        RECT  3.500 4.640 6.340 5.440 ;
        RECT  3.160 4.140 3.500 5.440 ;
        RECT  1.320 4.640 3.160 5.440 ;
        RECT  1.280 4.190 1.320 5.440 ;
        RECT  0.940 4.020 1.280 5.440 ;
        RECT  0.900 4.190 0.940 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.990 2.260 18.570 2.600 ;
        RECT  17.760 1.675 17.990 2.600 ;
        RECT  16.795 1.675 17.760 1.905 ;
        RECT  17.030 2.195 17.370 2.570 ;
        RECT  16.330 2.195 17.030 2.425 ;
        RECT  16.565 0.865 16.795 1.905 ;
        RECT  14.945 0.865 16.565 1.095 ;
        RECT  16.090 3.520 16.430 3.860 ;
        RECT  15.990 1.480 16.330 2.425 ;
        RECT  15.325 3.520 16.090 3.750 ;
        RECT  15.590 2.195 15.990 2.425 ;
        RECT  15.325 2.170 15.590 2.510 ;
        RECT  15.250 2.170 15.325 4.175 ;
        RECT  14.930 1.410 15.270 1.750 ;
        RECT  15.095 2.280 15.250 4.175 ;
        RECT  13.065 3.945 15.095 4.175 ;
        RECT  14.590 0.865 14.945 1.145 ;
        RECT  14.495 1.465 14.930 1.695 ;
        RECT  13.040 0.865 14.590 1.095 ;
        RECT  14.495 3.090 14.550 3.430 ;
        RECT  14.265 1.465 14.495 3.430 ;
        RECT  14.210 2.540 14.265 3.430 ;
        RECT  13.930 2.540 14.210 2.880 ;
        RECT  13.265 1.510 13.320 1.850 ;
        RECT  13.170 1.510 13.265 2.890 ;
        RECT  13.035 1.510 13.170 3.000 ;
        RECT  12.835 3.945 13.065 4.365 ;
        RECT  12.695 0.715 13.040 1.095 ;
        RECT  12.980 1.510 13.035 1.850 ;
        RECT  12.830 2.660 13.035 3.000 ;
        RECT  11.105 4.135 12.835 4.365 ;
        RECT  12.605 3.340 12.800 3.680 ;
        RECT  12.025 0.865 12.695 1.095 ;
        RECT  12.585 1.420 12.660 1.760 ;
        RECT  12.585 3.340 12.605 3.845 ;
        RECT  12.355 1.420 12.585 3.845 ;
        RECT  12.320 1.420 12.355 1.760 ;
        RECT  11.565 3.615 12.355 3.845 ;
        RECT  11.795 0.865 12.025 3.300 ;
        RECT  11.645 0.865 11.795 1.760 ;
        RECT  11.360 3.430 11.565 3.845 ;
        RECT  11.335 3.375 11.360 3.845 ;
        RECT  11.300 3.375 11.335 3.715 ;
        RECT  11.205 1.520 11.300 3.715 ;
        RECT  11.070 1.010 11.205 3.715 ;
        RECT  10.875 3.945 11.105 4.365 ;
        RECT  10.865 1.010 11.070 1.750 ;
        RECT  11.020 3.375 11.070 3.715 ;
        RECT  9.980 3.430 11.020 3.660 ;
        RECT  8.315 3.945 10.875 4.175 ;
        RECT  9.710 1.520 10.865 1.750 ;
        RECT  10.610 1.980 10.840 3.135 ;
        RECT  9.245 1.980 10.610 2.210 ;
        RECT  9.280 2.905 10.610 3.135 ;
        RECT  8.785 2.445 10.220 2.675 ;
        RECT  9.640 3.370 9.980 3.710 ;
        RECT  9.480 1.060 9.710 1.750 ;
        RECT  9.050 2.905 9.280 3.480 ;
        RECT  9.015 1.340 9.245 2.210 ;
        RECT  8.940 3.140 9.050 3.480 ;
        RECT  8.895 1.340 9.015 1.570 ;
        RECT  8.785 1.230 8.895 1.570 ;
        RECT  8.555 0.740 8.785 1.570 ;
        RECT  8.555 2.005 8.785 2.675 ;
        RECT  7.240 0.740 8.555 0.970 ;
        RECT  7.525 2.005 8.555 2.235 ;
        RECT  8.085 2.550 8.315 4.175 ;
        RECT  7.295 2.005 7.525 3.680 ;
        RECT  7.290 2.005 7.295 2.235 ;
        RECT  7.055 3.340 7.295 3.680 ;
        RECT  6.950 1.670 7.290 2.235 ;
        RECT  6.900 0.630 7.240 0.970 ;
        RECT  6.635 2.550 6.975 2.945 ;
        RECT  6.305 2.005 6.950 2.235 ;
        RECT  5.535 2.715 6.635 2.945 ;
        RECT  6.075 2.005 6.305 2.480 ;
        RECT  5.965 2.140 6.075 2.480 ;
        RECT  5.690 3.790 5.745 4.130 ;
        RECT  5.405 3.785 5.690 4.130 ;
        RECT  5.305 0.740 5.535 3.325 ;
        RECT  4.945 3.785 5.405 4.015 ;
        RECT  5.225 0.740 5.305 0.970 ;
        RECT  5.175 2.930 5.305 3.325 ;
        RECT  4.885 0.630 5.225 0.970 ;
        RECT  4.945 1.870 4.955 2.645 ;
        RECT  4.725 1.870 4.945 4.015 ;
        RECT  4.715 2.415 4.725 4.015 ;
        RECT  2.280 3.075 4.715 3.305 ;
        RECT  4.180 0.850 4.520 1.190 ;
        RECT  4.255 3.595 4.485 4.180 ;
        RECT  2.875 3.595 4.255 3.825 ;
        RECT  2.075 0.865 4.180 1.095 ;
        RECT  3.245 1.360 3.430 1.700 ;
        RECT  2.375 1.355 3.245 1.700 ;
        RECT  2.645 3.595 2.875 4.170 ;
        RECT  2.340 3.940 2.645 4.170 ;
        RECT  2.375 2.500 2.620 2.840 ;
        RECT  2.280 1.355 2.375 2.840 ;
        RECT  2.000 3.940 2.340 4.280 ;
        RECT  2.100 1.355 2.280 2.785 ;
        RECT  2.050 3.075 2.280 3.605 ;
        RECT  1.785 2.555 2.100 2.785 ;
        RECT  1.845 0.695 2.075 1.095 ;
        RECT  0.520 3.375 2.050 3.605 ;
        RECT  1.440 0.695 1.845 0.925 ;
        RECT  1.555 2.555 1.785 3.140 ;
        RECT  0.465 1.335 0.520 1.675 ;
        RECT  0.370 2.820 0.520 3.630 ;
        RECT  0.370 1.335 0.465 1.890 ;
        RECT  0.180 1.335 0.370 3.630 ;
        RECT  0.140 1.660 0.180 3.050 ;
    END
END SDFFRHQX2

MACRO SDFFRHQX1
    CLASS CORE ;
    FOREIGN SDFFRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRHQXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.290 2.380 3.745 2.635 ;
        RECT  3.005 2.050 3.290 2.635 ;
        RECT  2.950 2.050 3.005 2.390 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 1.460 1.845 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.250 2.910 15.040 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 1.245 16.335 3.195 ;
        RECT  16.270 1.245 16.330 4.085 ;
        RECT  16.105 1.245 16.270 4.290 ;
        RECT  15.210 1.245 16.105 1.475 ;
        RECT  16.055 2.965 16.105 4.290 ;
        RECT  15.930 3.480 16.055 4.290 ;
        RECT  14.980 0.730 15.210 1.475 ;
        RECT  14.870 0.730 14.980 1.070 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 1.750 4.480 2.110 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.170 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.930 -0.400 16.500 0.400 ;
        RECT  15.590 -0.400 15.930 0.950 ;
        RECT  14.445 -0.400 15.590 0.400 ;
        RECT  13.505 -0.400 14.445 0.575 ;
        RECT  12.365 -0.400 13.505 0.400 ;
        RECT  12.025 -0.400 12.365 0.575 ;
        RECT  9.435 -0.400 12.025 0.400 ;
        RECT  9.095 -0.400 9.435 1.130 ;
        RECT  6.660 -0.400 9.095 0.400 ;
        RECT  8.000 1.480 8.110 1.820 ;
        RECT  7.770 1.205 8.000 1.820 ;
        RECT  6.660 1.205 7.770 1.435 ;
        RECT  6.320 -0.400 6.660 1.435 ;
        RECT  3.140 -0.400 6.320 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.080 -0.400 2.800 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.990 4.640 16.500 5.440 ;
        RECT  14.650 3.535 14.990 5.440 ;
        RECT  14.010 3.535 14.650 3.765 ;
        RECT  12.730 4.640 14.650 5.440 ;
        RECT  13.920 2.985 14.010 3.765 ;
        RECT  13.780 2.930 13.920 3.765 ;
        RECT  13.580 2.930 13.780 3.270 ;
        RECT  12.315 4.465 12.730 5.440 ;
        RECT  9.855 4.640 12.315 5.440 ;
        RECT  9.440 4.465 9.855 5.440 ;
        RECT  6.680 4.640 9.440 5.440 ;
        RECT  6.340 3.980 6.680 5.440 ;
        RECT  3.500 4.640 6.340 5.440 ;
        RECT  3.160 4.140 3.500 5.440 ;
        RECT  0.920 4.640 3.160 5.440 ;
        RECT  0.580 3.850 0.920 5.440 ;
        RECT  0.000 4.640 0.580 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.350 1.710 15.690 2.050 ;
        RECT  14.400 1.710 15.350 1.940 ;
        RECT  13.795 2.450 15.330 2.680 ;
        RECT  14.170 0.865 14.400 1.940 ;
        RECT  13.925 4.000 14.265 4.340 ;
        RECT  12.725 0.865 14.170 1.095 ;
        RECT  13.345 4.000 13.925 4.285 ;
        RECT  13.795 1.375 13.845 1.715 ;
        RECT  13.565 1.375 13.795 2.680 ;
        RECT  13.505 1.375 13.565 1.715 ;
        RECT  13.345 2.210 13.565 2.680 ;
        RECT  13.225 2.210 13.345 4.285 ;
        RECT  13.115 2.405 13.225 4.285 ;
        RECT  8.425 3.945 13.115 4.175 ;
        RECT  12.705 1.410 13.045 1.750 ;
        RECT  12.355 0.865 12.725 1.145 ;
        RECT  12.600 1.520 12.705 1.750 ;
        RECT  12.370 1.520 12.600 3.500 ;
        RECT  12.260 2.580 12.370 3.500 ;
        RECT  11.780 0.865 12.355 1.095 ;
        RECT  12.040 2.580 12.260 2.920 ;
        RECT  11.550 0.865 11.780 3.600 ;
        RECT  11.000 0.865 11.550 1.105 ;
        RECT  11.310 3.370 11.550 3.600 ;
        RECT  11.120 1.605 11.315 1.945 ;
        RECT  10.970 3.370 11.310 3.710 ;
        RECT  10.975 1.605 11.120 3.055 ;
        RECT  10.715 0.865 11.000 1.275 ;
        RECT  10.890 1.660 10.975 3.055 ;
        RECT  10.660 0.935 10.715 1.275 ;
        RECT  10.430 1.595 10.660 3.710 ;
        RECT  10.425 1.595 10.430 1.825 ;
        RECT  10.250 3.370 10.430 3.710 ;
        RECT  10.200 1.120 10.425 1.825 ;
        RECT  10.195 1.010 10.200 1.825 ;
        RECT  9.965 2.300 10.200 2.705 ;
        RECT  9.860 1.010 10.195 1.350 ;
        RECT  9.735 1.640 9.965 3.580 ;
        RECT  8.940 1.640 9.735 1.870 ;
        RECT  9.270 3.350 9.735 3.580 ;
        RECT  9.275 2.105 9.505 2.915 ;
        RECT  7.450 2.105 9.275 2.335 ;
        RECT  8.930 3.350 9.270 3.690 ;
        RECT  8.805 1.530 8.940 1.870 ;
        RECT  8.575 0.685 8.805 1.870 ;
        RECT  6.960 0.685 8.575 0.915 ;
        RECT  8.300 2.635 8.425 4.175 ;
        RECT  8.195 2.580 8.300 4.175 ;
        RECT  7.960 2.580 8.195 2.920 ;
        RECT  7.310 1.725 7.450 3.680 ;
        RECT  7.220 1.670 7.310 3.680 ;
        RECT  6.970 1.670 7.220 2.010 ;
        RECT  7.050 3.340 7.220 3.680 ;
        RECT  6.760 2.580 6.990 2.945 ;
        RECT  6.270 1.780 6.970 2.010 ;
        RECT  5.535 2.715 6.760 2.945 ;
        RECT  6.040 1.780 6.270 2.370 ;
        RECT  5.930 2.030 6.040 2.370 ;
        RECT  5.470 3.740 5.810 4.080 ;
        RECT  5.435 1.045 5.535 2.945 ;
        RECT  4.945 3.740 5.470 3.970 ;
        RECT  5.305 1.045 5.435 3.325 ;
        RECT  5.300 1.045 5.305 1.275 ;
        RECT  5.205 2.715 5.305 3.325 ;
        RECT  4.960 0.935 5.300 1.275 ;
        RECT  4.715 1.830 4.945 3.970 ;
        RECT  2.300 3.075 4.715 3.305 ;
        RECT  4.160 0.865 4.500 1.230 ;
        RECT  4.255 3.595 4.485 4.040 ;
        RECT  2.760 3.595 4.255 3.825 ;
        RECT  1.780 0.865 4.160 1.095 ;
        RECT  3.415 1.330 3.420 1.670 ;
        RECT  3.080 1.330 3.415 1.690 ;
        RECT  2.435 1.460 3.080 1.690 ;
        RECT  2.530 3.595 2.760 4.170 ;
        RECT  2.435 2.500 2.590 2.840 ;
        RECT  2.340 3.940 2.530 4.170 ;
        RECT  2.250 1.460 2.435 2.840 ;
        RECT  2.000 3.940 2.340 4.280 ;
        RECT  2.070 3.075 2.300 3.610 ;
        RECT  2.145 1.460 2.250 2.785 ;
        RECT  2.090 1.460 2.145 1.800 ;
        RECT  1.840 2.555 2.145 2.785 ;
        RECT  0.520 3.380 2.070 3.610 ;
        RECT  1.610 2.555 1.840 3.140 ;
        RECT  1.440 0.640 1.780 1.095 ;
        RECT  1.500 2.800 1.610 3.140 ;
        RECT  0.395 1.330 0.520 1.670 ;
        RECT  0.395 2.890 0.520 3.610 ;
        RECT  0.290 1.330 0.395 3.610 ;
        RECT  0.165 1.330 0.290 3.230 ;
    END
END SDFFRHQX1

MACRO SDFFRXL
    CLASS CORE ;
    FOREIGN SDFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 2.320 3.790 2.675 ;
        RECT  3.335 2.320 3.675 2.925 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 1.800 1.810 2.290 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.270 2.900 7.610 3.240 ;
        RECT  7.120 2.900 7.270 3.220 ;
        RECT  7.045 2.360 7.120 3.220 ;
        RECT  6.890 2.360 7.045 3.185 ;
        RECT  6.760 2.360 6.890 2.680 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.765 0.865 16.995 4.035 ;
        RECT  16.410 0.865 16.765 1.095 ;
        RECT  16.615 3.500 16.765 4.035 ;
        RECT  16.490 3.805 16.615 4.035 ;
        RECT  16.150 3.805 16.490 4.230 ;
        RECT  16.070 0.635 16.410 1.095 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.135 3.620 18.220 3.960 ;
        RECT  17.905 1.890 18.135 3.960 ;
        RECT  17.820 1.890 17.905 2.120 ;
        RECT  17.880 3.620 17.905 3.960 ;
        RECT  17.300 1.190 17.820 2.120 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.105 1.575 4.495 2.105 ;
        RECT  4.035 1.715 4.105 2.080 ;
        RECT  3.980 1.740 4.035 2.080 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.715 1.180 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.140 -0.400 18.480 0.400 ;
        RECT  16.800 -0.400 17.140 0.575 ;
        RECT  15.530 -0.400 16.800 0.400 ;
        RECT  15.190 -0.400 15.530 0.950 ;
        RECT  13.770 -0.400 15.190 0.400 ;
        RECT  13.430 -0.400 13.770 1.110 ;
        RECT  9.005 -0.400 13.430 0.400 ;
        RECT  10.535 1.205 10.875 1.760 ;
        RECT  9.300 1.205 10.535 1.435 ;
        RECT  9.005 1.205 9.300 1.580 ;
        RECT  8.960 -0.400 9.005 1.580 ;
        RECT  8.775 -0.400 8.960 1.525 ;
        RECT  6.990 -0.400 8.775 0.400 ;
        RECT  6.650 -0.400 6.990 0.960 ;
        RECT  3.300 -0.400 6.650 0.400 ;
        RECT  2.960 -0.400 3.300 0.575 ;
        RECT  1.210 -0.400 2.960 0.400 ;
        RECT  0.870 -0.400 1.210 0.575 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.450 4.640 18.480 5.440 ;
        RECT  17.110 4.465 17.450 5.440 ;
        RECT  15.730 4.640 17.110 5.440 ;
        RECT  15.390 4.090 15.730 5.440 ;
        RECT  13.705 4.640 15.390 5.440 ;
        RECT  13.365 4.080 13.705 5.440 ;
        RECT  11.370 4.640 13.365 5.440 ;
        RECT  10.430 4.080 11.370 5.440 ;
        RECT  7.370 4.640 10.430 5.440 ;
        RECT  7.030 4.465 7.370 5.440 ;
        RECT  3.730 4.640 7.030 5.440 ;
        RECT  3.390 4.080 3.730 5.440 ;
        RECT  0.760 4.640 3.390 5.440 ;
        RECT  0.420 4.465 0.760 5.440 ;
        RECT  0.000 4.640 0.420 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.380 1.380 16.490 3.160 ;
        RECT  16.150 1.380 16.380 3.350 ;
        RECT  15.970 1.380 16.150 1.850 ;
        RECT  16.040 2.820 16.150 3.350 ;
        RECT  15.625 1.880 15.670 2.220 ;
        RECT  15.615 1.865 15.625 2.220 ;
        RECT  15.115 1.865 15.615 2.245 ;
        RECT  14.885 1.865 15.115 3.850 ;
        RECT  14.675 1.865 14.885 2.095 ;
        RECT  14.410 3.620 14.885 3.850 ;
        RECT  14.445 0.915 14.675 2.095 ;
        RECT  14.310 3.005 14.650 3.390 ;
        RECT  14.285 0.915 14.445 1.825 ;
        RECT  14.070 3.620 14.410 3.960 ;
        RECT  13.175 3.160 14.310 3.390 ;
        RECT  13.930 1.595 14.285 1.825 ;
        RECT  13.700 1.595 13.930 2.580 ;
        RECT  13.590 2.240 13.700 2.580 ;
        RECT  12.995 1.400 13.175 3.405 ;
        RECT  12.995 4.000 13.000 4.340 ;
        RECT  12.945 1.400 12.995 4.340 ;
        RECT  12.230 1.400 12.945 1.630 ;
        RECT  12.765 3.160 12.945 4.340 ;
        RECT  12.660 4.000 12.765 4.340 ;
        RECT  12.540 2.390 12.595 2.730 ;
        RECT  12.255 2.390 12.540 2.875 ;
        RECT  12.175 2.645 12.255 2.875 ;
        RECT  11.890 1.290 12.230 1.630 ;
        RECT  11.945 2.645 12.175 3.850 ;
        RECT  10.495 3.620 11.945 3.850 ;
        RECT  11.575 2.035 11.880 2.375 ;
        RECT  11.345 0.675 11.575 3.385 ;
        RECT  9.670 0.675 11.345 0.905 ;
        RECT  10.730 3.155 11.345 3.385 ;
        RECT  9.615 2.140 11.030 2.480 ;
        RECT  10.265 2.810 10.495 3.850 ;
        RECT  10.135 3.620 10.265 3.850 ;
        RECT  9.905 3.620 10.135 4.365 ;
        RECT  7.830 4.135 9.905 4.365 ;
        RECT  9.330 0.635 9.670 0.975 ;
        RECT  9.385 1.825 9.615 3.690 ;
        RECT  8.435 1.825 9.385 2.055 ;
        RECT  9.080 3.460 9.385 3.690 ;
        RECT  8.740 3.460 9.080 3.800 ;
        RECT  8.730 2.440 9.070 2.780 ;
        RECT  8.290 2.495 8.730 2.725 ;
        RECT  8.205 1.100 8.435 2.055 ;
        RECT  8.060 2.435 8.290 3.870 ;
        RECT  8.095 1.100 8.205 1.885 ;
        RECT  6.540 1.655 8.095 1.885 ;
        RECT  7.895 2.435 8.060 2.665 ;
        RECT  7.555 2.115 7.895 2.665 ;
        RECT  7.600 4.005 7.830 4.365 ;
        RECT  7.535 0.770 7.805 1.110 ;
        RECT  6.645 4.005 7.600 4.235 ;
        RECT  7.465 0.770 7.535 1.420 ;
        RECT  7.305 0.825 7.465 1.420 ;
        RECT  5.935 1.190 7.305 1.420 ;
        RECT  6.495 4.005 6.645 4.355 ;
        RECT  6.200 1.655 6.540 2.080 ;
        RECT  6.415 4.005 6.495 4.410 ;
        RECT  6.155 4.070 6.415 4.410 ;
        RECT  5.625 4.125 6.155 4.355 ;
        RECT  5.935 2.505 6.085 3.800 ;
        RECT  5.855 1.190 5.935 3.800 ;
        RECT  5.705 1.190 5.855 2.735 ;
        RECT  5.500 1.190 5.705 1.420 ;
        RECT  5.395 2.970 5.625 4.355 ;
        RECT  5.160 0.980 5.500 1.420 ;
        RECT  5.200 2.970 5.395 3.200 ;
        RECT  4.275 4.125 5.395 4.355 ;
        RECT  5.090 1.945 5.200 3.200 ;
        RECT  4.935 3.460 5.165 3.800 ;
        RECT  4.970 1.890 5.090 3.200 ;
        RECT  4.750 1.890 4.970 2.230 ;
        RECT  4.740 3.460 4.935 3.690 ;
        RECT  4.510 3.160 4.740 3.690 ;
        RECT  4.570 0.960 4.660 1.300 ;
        RECT  4.320 0.865 4.570 1.300 ;
        RECT  2.710 3.160 4.510 3.390 ;
        RECT  2.155 0.865 4.320 1.095 ;
        RECT  4.045 3.620 4.275 4.355 ;
        RECT  3.155 3.620 4.045 3.850 ;
        RECT  3.170 1.615 3.510 1.955 ;
        RECT  2.430 1.670 3.170 1.900 ;
        RECT  2.925 3.620 3.155 4.225 ;
        RECT  1.395 3.995 2.925 4.225 ;
        RECT  2.370 3.050 2.710 3.390 ;
        RECT  2.375 1.450 2.430 1.900 ;
        RECT  2.375 2.480 2.380 2.820 ;
        RECT  2.145 1.450 2.375 2.820 ;
        RECT  1.940 0.685 2.155 1.095 ;
        RECT  2.090 1.450 2.145 1.790 ;
        RECT  2.040 2.480 2.145 2.820 ;
        RECT  1.935 2.590 2.040 2.820 ;
        RECT  1.935 3.425 1.990 3.765 ;
        RECT  1.925 0.630 1.940 1.095 ;
        RECT  1.705 2.590 1.935 3.765 ;
        RECT  1.600 0.630 1.925 0.970 ;
        RECT  1.650 3.425 1.705 3.765 ;
        RECT  1.165 3.745 1.395 4.225 ;
        RECT  0.540 3.745 1.165 3.975 ;
        RECT  0.395 1.230 0.540 1.570 ;
        RECT  0.395 3.530 0.540 3.975 ;
        RECT  0.165 1.230 0.395 3.975 ;
    END
END SDFFRXL

MACRO SDFFRX4
    CLASS CORE ;
    FOREIGN SDFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 2.050 3.165 2.785 ;
        RECT  2.780 2.060 2.825 2.785 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.290 1.780 2.340 ;
        RECT  1.470 1.285 1.765 2.340 ;
        RECT  1.430 1.285 1.470 2.300 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.320 2.745 7.780 3.495 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.600 1.195 20.980 3.220 ;
        RECT  20.580 1.195 20.600 1.535 ;
        RECT  20.580 2.780 20.600 3.120 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.200 1.260 22.300 3.120 ;
        RECT  21.920 1.195 22.200 3.120 ;
        RECT  21.915 1.195 21.920 2.075 ;
        RECT  21.860 2.780 21.920 3.120 ;
        RECT  21.860 1.195 21.915 1.535 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.945 2.360 4.175 2.700 ;
        RECT  3.815 2.360 3.945 2.590 ;
        RECT  3.585 1.845 3.815 2.590 ;
        RECT  3.515 1.845 3.585 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.660 2.350 1.120 2.835 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.840 -0.400 23.100 0.400 ;
        RECT  22.500 -0.400 22.840 0.950 ;
        RECT  21.560 -0.400 22.500 0.400 ;
        RECT  21.220 -0.400 21.560 0.950 ;
        RECT  20.280 -0.400 21.220 0.400 ;
        RECT  19.940 -0.400 20.280 0.950 ;
        RECT  18.910 -0.400 19.940 0.400 ;
        RECT  18.570 -0.400 18.910 0.950 ;
        RECT  17.470 -0.400 18.570 0.400 ;
        RECT  17.130 -0.400 17.470 0.950 ;
        RECT  16.010 -0.400 17.130 0.400 ;
        RECT  15.670 -0.400 16.010 0.950 ;
        RECT  14.240 -0.400 15.670 0.400 ;
        RECT  13.900 -0.400 14.240 1.080 ;
        RECT  11.645 -0.400 13.900 0.400 ;
        RECT  11.415 -0.400 11.645 1.475 ;
        RECT  9.790 -0.400 11.415 0.400 ;
        RECT  11.270 1.245 11.415 1.475 ;
        RECT  9.450 -0.400 9.790 0.960 ;
        RECT  7.780 -0.400 9.450 0.400 ;
        RECT  7.440 -0.400 7.780 1.335 ;
        RECT  3.240 -0.400 7.440 0.400 ;
        RECT  2.900 -0.400 3.240 0.575 ;
        RECT  1.080 -0.400 2.900 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.840 4.640 23.100 5.440 ;
        RECT  22.500 4.040 22.840 5.440 ;
        RECT  21.560 4.640 22.500 5.440 ;
        RECT  21.220 4.040 21.560 5.440 ;
        RECT  20.280 4.640 21.220 5.440 ;
        RECT  19.940 4.080 20.280 5.440 ;
        RECT  18.710 4.640 19.940 5.440 ;
        RECT  18.370 3.055 18.710 5.440 ;
        RECT  16.110 4.640 18.370 5.440 ;
        RECT  15.770 4.080 16.110 5.440 ;
        RECT  13.630 4.640 15.770 5.440 ;
        RECT  13.290 3.675 13.630 5.440 ;
        RECT  10.780 4.640 13.290 5.440 ;
        RECT  10.440 3.920 10.780 5.440 ;
        RECT  7.120 4.640 10.440 5.440 ;
        RECT  6.780 4.465 7.120 5.440 ;
        RECT  3.880 4.640 6.780 5.440 ;
        RECT  3.540 4.080 3.880 5.440 ;
        RECT  0.850 4.640 3.540 5.440 ;
        RECT  0.510 4.465 0.850 5.440 ;
        RECT  0.000 4.640 0.510 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.605 2.030 22.835 3.750 ;
        RECT  20.275 3.520 22.605 3.750 ;
        RECT  20.045 1.395 20.275 3.750 ;
        RECT  19.590 1.395 20.045 1.730 ;
        RECT  19.430 3.265 20.045 3.495 ;
        RECT  18.810 2.100 19.750 2.440 ;
        RECT  19.250 1.390 19.590 1.730 ;
        RECT  19.090 2.975 19.430 3.785 ;
        RECT  19.240 1.395 19.250 1.675 ;
        RECT  18.190 2.155 18.810 2.385 ;
        RECT  17.960 0.720 18.190 2.690 ;
        RECT  17.850 0.720 17.960 1.475 ;
        RECT  17.430 2.460 17.960 2.690 ;
        RECT  16.750 1.245 17.850 1.475 ;
        RECT  17.355 1.725 17.710 2.065 ;
        RECT  17.200 2.460 17.430 3.835 ;
        RECT  16.770 1.725 17.355 2.105 ;
        RECT  17.090 2.985 17.200 3.835 ;
        RECT  15.500 3.605 17.090 3.835 ;
        RECT  15.765 1.875 16.770 2.105 ;
        RECT  16.520 0.700 16.750 1.475 ;
        RECT  16.410 0.700 16.520 1.040 ;
        RECT  15.535 1.495 15.765 3.365 ;
        RECT  13.195 1.495 15.535 1.735 ;
        RECT  14.905 3.135 15.535 3.365 ;
        RECT  15.270 3.605 15.500 4.250 ;
        RECT  14.765 2.425 15.105 2.820 ;
        RECT  14.905 3.750 14.960 4.090 ;
        RECT  14.675 3.135 14.905 4.090 ;
        RECT  12.735 2.425 14.765 2.655 ;
        RECT  12.995 3.135 14.675 3.365 ;
        RECT  14.620 3.750 14.675 4.090 ;
        RECT  12.965 1.095 13.195 1.735 ;
        RECT  12.765 3.135 12.995 3.855 ;
        RECT  12.550 1.095 12.965 1.325 ;
        RECT  12.350 3.625 12.765 3.855 ;
        RECT  12.505 1.740 12.735 2.655 ;
        RECT  12.220 2.425 12.505 2.655 ;
        RECT  12.010 3.625 12.350 3.990 ;
        RECT  11.990 1.745 12.220 3.145 ;
        RECT  10.765 1.745 11.990 1.975 ;
        RECT  11.545 2.915 11.990 3.145 ;
        RECT  10.175 2.230 11.760 2.460 ;
        RECT  11.540 2.915 11.545 3.945 ;
        RECT  11.315 2.915 11.540 4.000 ;
        RECT  11.200 3.660 11.315 4.000 ;
        RECT  10.805 2.840 10.970 3.180 ;
        RECT  10.575 2.840 10.805 3.660 ;
        RECT  10.535 0.675 10.765 1.975 ;
        RECT  10.045 3.430 10.575 3.660 ;
        RECT  10.040 0.675 10.535 0.905 ;
        RECT  9.945 1.565 10.175 3.145 ;
        RECT  9.815 3.430 10.045 4.365 ;
        RECT  9.230 1.565 9.945 1.795 ;
        RECT  9.500 2.915 9.945 3.145 ;
        RECT  7.665 4.135 9.815 4.365 ;
        RECT  9.160 2.915 9.500 3.870 ;
        RECT  9.130 2.100 9.470 2.440 ;
        RECT  8.890 1.430 9.230 1.795 ;
        RECT  8.315 2.155 9.130 2.385 ;
        RECT  6.960 1.565 8.890 1.795 ;
        RECT  8.315 3.560 8.370 3.900 ;
        RECT  8.085 2.025 8.315 3.900 ;
        RECT  7.570 2.025 8.085 2.255 ;
        RECT  8.030 3.560 8.085 3.900 ;
        RECT  7.435 3.945 7.665 4.365 ;
        RECT  6.465 3.945 7.435 4.175 ;
        RECT  6.730 1.565 6.960 2.660 ;
        RECT  5.625 0.825 6.950 1.055 ;
        RECT  6.620 2.320 6.730 2.660 ;
        RECT  6.310 3.035 6.465 4.345 ;
        RECT  6.235 1.980 6.310 4.345 ;
        RECT  6.080 1.980 6.235 3.265 ;
        RECT  4.365 4.115 6.235 4.345 ;
        RECT  5.095 1.980 6.080 2.210 ;
        RECT  5.665 3.500 5.920 3.840 ;
        RECT  5.435 2.465 5.665 3.840 ;
        RECT  5.400 0.825 5.625 1.415 ;
        RECT  4.635 2.465 5.435 2.695 ;
        RECT  5.395 0.825 5.400 1.470 ;
        RECT  5.345 1.130 5.395 1.470 ;
        RECT  5.060 1.130 5.345 1.635 ;
        RECT  5.025 3.430 5.200 3.770 ;
        RECT  4.865 1.870 5.095 2.210 ;
        RECT  4.635 1.405 5.060 1.635 ;
        RECT  4.795 3.135 5.025 3.770 ;
        RECT  2.760 3.135 4.795 3.365 ;
        RECT  4.405 1.405 4.635 2.695 ;
        RECT  4.260 0.830 4.600 1.170 ;
        RECT  4.135 3.615 4.365 4.345 ;
        RECT  2.615 0.865 4.260 1.095 ;
        RECT  3.240 3.615 4.135 3.845 ;
        RECT  2.475 1.345 3.520 1.575 ;
        RECT  3.010 3.615 3.240 4.235 ;
        RECT  0.520 4.005 3.010 4.235 ;
        RECT  2.475 3.135 2.760 3.600 ;
        RECT  2.385 0.680 2.615 1.095 ;
        RECT  2.145 1.345 2.475 2.845 ;
        RECT  2.420 3.260 2.475 3.600 ;
        RECT  1.540 0.680 2.385 0.910 ;
        RECT  2.070 1.360 2.145 1.700 ;
        RECT  2.105 2.615 2.145 2.845 ;
        RECT  1.875 2.615 2.105 3.650 ;
        RECT  1.840 3.420 1.875 3.650 ;
        RECT  1.500 3.420 1.840 3.760 ;
        RECT  0.405 1.265 0.520 1.605 ;
        RECT  0.405 3.180 0.520 4.235 ;
        RECT  0.290 1.265 0.405 4.235 ;
        RECT  0.175 1.265 0.290 3.520 ;
    END
END SDFFRX4

MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.830 2.260 3.435 2.680 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.240 1.795 1.560 ;
        RECT  1.715 1.930 1.770 2.270 ;
        RECT  1.485 1.240 1.715 2.270 ;
        RECT  1.430 1.930 1.485 2.270 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.245 2.875 7.300 3.390 ;
        RECT  6.960 2.755 7.245 3.390 ;
        RECT  6.815 2.755 6.960 3.335 ;
        RECT  6.770 2.875 6.815 3.240 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.205 1.825 18.265 2.075 ;
        RECT  18.205 2.930 18.260 3.270 ;
        RECT  18.020 1.825 18.205 3.270 ;
        RECT  17.975 1.370 18.020 3.270 ;
        RECT  17.790 1.370 17.975 2.055 ;
        RECT  17.920 2.930 17.975 3.270 ;
        RECT  17.680 1.370 17.790 1.710 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.580 0.955 19.645 3.230 ;
        RECT  19.570 0.955 19.580 3.270 ;
        RECT  19.345 0.685 19.570 3.270 ;
        RECT  19.230 0.685 19.345 1.625 ;
        RECT  19.240 2.910 19.345 3.270 ;
        RECT  19.210 2.930 19.240 3.270 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.840 1.550 4.480 2.120 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.965 1.800 1.150 2.120 ;
        RECT  0.625 1.715 0.965 2.820 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.735 -0.400 19.800 0.400 ;
        RECT  18.505 -0.400 18.735 1.555 ;
        RECT  16.760 -0.400 18.505 0.400 ;
        RECT  16.420 -0.400 16.760 1.190 ;
        RECT  15.270 -0.400 16.420 0.400 ;
        RECT  14.930 -0.400 15.270 0.575 ;
        RECT  13.410 -0.400 14.930 0.400 ;
        RECT  13.070 -0.400 13.410 1.250 ;
        RECT  10.680 -0.400 13.070 0.400 ;
        RECT  10.340 -0.400 10.680 1.370 ;
        RECT  8.980 -0.400 10.340 0.400 ;
        RECT  8.640 -0.400 8.980 0.960 ;
        RECT  7.760 -0.400 8.640 0.440 ;
        RECT  7.335 -0.400 7.760 1.335 ;
        RECT  3.140 -0.400 7.335 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.080 -0.400 2.800 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.900 4.640 19.800 5.440 ;
        RECT  18.560 4.080 18.900 5.440 ;
        RECT  16.840 4.640 18.560 5.440 ;
        RECT  16.500 3.680 16.840 5.440 ;
        RECT  14.060 4.640 16.500 5.440 ;
        RECT  13.720 4.080 14.060 5.440 ;
        RECT  11.345 4.640 13.720 5.440 ;
        RECT  9.900 4.135 11.345 5.440 ;
        RECT  7.000 4.640 9.900 5.440 ;
        RECT  6.660 4.465 7.000 5.440 ;
        RECT  3.840 4.640 6.660 5.440 ;
        RECT  3.500 3.980 3.840 5.440 ;
        RECT  1.080 4.640 3.500 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.885 1.910 19.115 2.655 ;
        RECT  18.840 2.425 18.885 2.655 ;
        RECT  18.610 2.425 18.840 3.805 ;
        RECT  17.560 3.575 18.610 3.805 ;
        RECT  17.450 3.575 17.560 4.020 ;
        RECT  17.450 0.665 17.520 1.005 ;
        RECT  17.220 0.665 17.450 4.020 ;
        RECT  17.180 0.665 17.220 1.005 ;
        RECT  16.935 1.590 16.990 2.045 ;
        RECT  16.705 1.590 16.935 3.165 ;
        RECT  16.650 1.590 16.705 2.045 ;
        RECT  16.160 2.935 16.705 3.165 ;
        RECT  16.040 1.815 16.650 2.045 ;
        RECT  15.930 2.935 16.160 3.510 ;
        RECT  15.810 0.910 16.040 2.045 ;
        RECT  15.380 3.280 15.930 3.510 ;
        RECT  15.700 0.910 15.810 1.250 ;
        RECT  15.130 1.815 15.810 2.045 ;
        RECT  15.270 3.280 15.380 3.620 ;
        RECT  15.040 3.280 15.270 4.270 ;
        RECT  14.690 2.460 15.190 2.800 ;
        RECT  14.845 1.630 15.130 2.045 ;
        RECT  14.760 3.930 15.040 4.270 ;
        RECT  14.790 1.630 14.845 1.970 ;
        RECT  14.560 2.460 14.690 3.335 ;
        RECT  14.330 1.685 14.560 3.335 ;
        RECT  14.230 1.685 14.330 1.915 ;
        RECT  14.320 2.680 14.330 3.335 ;
        RECT  13.305 3.105 14.320 3.335 ;
        RECT  14.000 1.225 14.230 1.915 ;
        RECT  14.045 2.205 14.100 2.435 ;
        RECT  13.815 2.205 14.045 2.440 ;
        RECT  13.770 1.225 14.000 1.755 ;
        RECT  13.425 2.210 13.815 2.440 ;
        RECT  12.100 1.525 13.770 1.755 ;
        RECT  13.195 1.985 13.425 2.440 ;
        RECT  13.075 3.105 13.305 3.480 ;
        RECT  11.640 1.985 13.195 2.215 ;
        RECT  12.740 3.250 13.075 3.480 ;
        RECT  12.400 3.250 12.740 3.590 ;
        RECT  12.160 2.600 12.500 2.940 ;
        RECT  12.145 2.710 12.160 2.940 ;
        RECT  11.915 2.710 12.145 3.900 ;
        RECT  11.870 1.090 12.100 1.755 ;
        RECT  10.015 3.670 11.915 3.900 ;
        RECT  11.700 1.090 11.870 1.430 ;
        RECT  11.410 1.705 11.640 3.435 ;
        RECT  9.880 1.705 11.410 1.935 ;
        RECT  10.470 3.205 11.410 3.435 ;
        RECT  10.840 2.170 11.180 2.885 ;
        RECT  9.215 2.170 10.840 2.400 ;
        RECT  10.170 2.630 10.510 2.970 ;
        RECT  10.015 2.685 10.170 2.970 ;
        RECT  9.785 2.685 10.015 3.900 ;
        RECT  9.875 1.205 9.880 1.935 ;
        RECT  9.765 1.150 9.875 1.935 ;
        RECT  9.575 3.670 9.785 3.900 ;
        RECT  9.590 0.665 9.765 1.935 ;
        RECT  9.535 0.665 9.590 1.490 ;
        RECT  9.345 3.670 9.575 4.355 ;
        RECT  9.270 0.665 9.535 0.895 ;
        RECT  7.465 4.125 9.345 4.355 ;
        RECT  8.985 1.575 9.215 3.185 ;
        RECT  8.480 1.575 8.985 1.805 ;
        RECT  8.795 2.955 8.985 3.185 ;
        RECT  8.795 3.470 8.850 3.810 ;
        RECT  8.565 2.955 8.795 3.810 ;
        RECT  8.415 2.140 8.755 2.480 ;
        RECT  8.510 3.470 8.565 3.810 ;
        RECT  8.250 1.455 8.480 1.805 ;
        RECT  7.985 2.195 8.415 2.425 ;
        RECT  8.140 1.455 8.250 1.795 ;
        RECT  6.320 1.565 8.140 1.795 ;
        RECT  7.985 3.550 8.040 3.890 ;
        RECT  7.755 2.195 7.985 3.890 ;
        RECT  7.750 2.195 7.755 2.425 ;
        RECT  7.700 3.550 7.755 3.890 ;
        RECT  7.200 2.030 7.750 2.425 ;
        RECT  7.235 3.945 7.465 4.355 ;
        RECT  6.345 3.945 7.235 4.175 ;
        RECT  6.720 0.675 7.060 1.110 ;
        RECT  5.665 0.675 6.720 0.905 ;
        RECT  6.115 3.945 6.345 4.255 ;
        RECT  5.990 1.565 6.320 2.085 ;
        RECT  5.200 4.025 6.115 4.255 ;
        RECT  5.980 1.745 5.990 2.085 ;
        RECT  5.685 3.300 5.740 3.640 ;
        RECT  5.665 3.280 5.685 3.640 ;
        RECT  5.435 0.675 5.665 3.640 ;
        RECT  4.960 0.930 5.435 1.270 ;
        RECT  5.400 3.300 5.435 3.640 ;
        RECT  5.100 3.970 5.200 4.310 ;
        RECT  5.055 1.655 5.100 4.310 ;
        RECT  4.870 1.600 5.055 4.310 ;
        RECT  4.715 1.600 4.870 1.940 ;
        RECT  4.860 3.970 4.870 4.310 ;
        RECT  4.385 3.970 4.860 4.200 ;
        RECT  4.205 2.850 4.545 3.190 ;
        RECT  4.160 0.865 4.500 1.270 ;
        RECT  4.155 3.450 4.385 4.200 ;
        RECT  2.475 2.935 4.205 3.165 ;
        RECT  2.565 0.865 4.160 1.095 ;
        RECT  2.515 3.450 4.155 3.680 ;
        RECT  3.020 1.635 3.360 1.975 ;
        RECT  2.410 1.690 3.020 1.920 ;
        RECT  2.335 0.665 2.565 1.095 ;
        RECT  2.285 3.450 2.515 4.235 ;
        RECT  2.230 1.460 2.410 2.070 ;
        RECT  1.785 0.665 2.335 0.895 ;
        RECT  0.520 4.005 2.285 4.235 ;
        RECT  2.070 1.460 2.230 2.740 ;
        RECT  2.065 1.840 2.070 2.740 ;
        RECT  2.000 1.840 2.065 3.180 ;
        RECT  1.880 2.505 2.000 3.180 ;
        RECT  1.835 2.505 1.880 3.770 ;
        RECT  1.650 2.840 1.835 3.770 ;
        RECT  1.440 0.665 1.785 0.960 ;
        RECT  1.540 3.430 1.650 3.770 ;
        RECT  0.395 1.100 0.520 1.440 ;
        RECT  0.395 3.630 0.520 4.235 ;
        RECT  0.165 1.100 0.395 4.235 ;
    END
END SDFFRX2

MACRO SDFFRX1
    CLASS CORE ;
    FOREIGN SDFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 2.520 3.710 2.860 ;
        RECT  3.370 2.400 3.620 2.860 ;
        RECT  3.360 2.400 3.370 2.820 ;
        RECT  3.130 2.400 3.360 2.660 ;
        RECT  2.840 2.390 3.130 2.660 ;
        RECT  2.780 2.390 2.840 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.760 1.810 2.220 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.165 3.340 7.795 3.570 ;
        RECT  6.935 2.390 7.165 3.570 ;
        RECT  6.770 2.390 6.935 2.650 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.150 2.035 17.380 3.295 ;
        RECT  16.715 2.035 17.150 2.265 ;
        RECT  17.020 3.065 17.150 3.295 ;
        RECT  16.715 3.065 17.020 3.790 ;
        RECT  16.585 1.820 16.715 2.265 ;
        RECT  16.490 3.525 16.715 3.790 ;
        RECT  16.355 1.380 16.585 2.265 ;
        RECT  16.150 3.525 16.490 3.990 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.965 1.355 17.980 1.695 ;
        RECT  17.750 1.270 17.965 3.930 ;
        RECT  17.705 1.270 17.750 3.980 ;
        RECT  17.640 1.270 17.705 1.695 ;
        RECT  17.410 3.640 17.705 3.980 ;
        RECT  17.375 1.270 17.640 1.655 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 1.730 4.320 2.100 ;
        RECT  3.440 1.820 3.980 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.670 1.180 3.230 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.210 -0.400 18.480 0.400 ;
        RECT  16.870 -0.400 17.210 0.575 ;
        RECT  15.215 -0.400 16.870 0.400 ;
        RECT  14.875 -0.400 15.215 0.575 ;
        RECT  13.660 -0.400 14.875 0.400 ;
        RECT  13.320 -0.400 13.660 1.310 ;
        RECT  9.005 -0.400 13.320 0.400 ;
        RECT  10.780 1.440 10.890 1.780 ;
        RECT  10.550 1.205 10.780 1.780 ;
        RECT  9.300 1.205 10.550 1.435 ;
        RECT  9.005 1.205 9.300 1.525 ;
        RECT  8.775 -0.400 9.005 1.525 ;
        RECT  6.990 -0.400 8.775 0.400 ;
        RECT  6.650 -0.400 6.990 0.960 ;
        RECT  3.200 -0.400 6.650 0.400 ;
        RECT  2.860 -0.400 3.200 0.575 ;
        RECT  0.585 -0.400 2.860 0.400 ;
        RECT  0.245 -0.400 0.585 0.575 ;
        RECT  0.000 -0.400 0.245 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.070 4.640 18.480 5.440 ;
        RECT  16.730 4.465 17.070 5.440 ;
        RECT  15.730 4.640 16.730 5.440 ;
        RECT  15.390 3.620 15.730 5.440 ;
        RECT  13.710 4.640 15.390 5.440 ;
        RECT  13.370 4.070 13.710 5.440 ;
        RECT  11.370 4.640 13.370 5.440 ;
        RECT  10.430 4.070 11.370 5.440 ;
        RECT  7.300 4.640 10.430 5.440 ;
        RECT  6.960 4.465 7.300 5.440 ;
        RECT  3.730 4.640 6.960 5.440 ;
        RECT  3.390 4.080 3.730 5.440 ;
        RECT  1.130 4.640 3.390 5.440 ;
        RECT  0.790 4.465 1.130 5.440 ;
        RECT  0.000 4.640 0.790 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.390 2.495 16.920 2.835 ;
        RECT  16.115 2.495 16.390 3.140 ;
        RECT  16.050 1.250 16.115 3.140 ;
        RECT  15.815 1.250 16.050 2.795 ;
        RECT  15.760 1.250 15.815 1.550 ;
        RECT  15.420 1.210 15.760 1.550 ;
        RECT  15.425 1.825 15.530 2.110 ;
        RECT  15.195 1.825 15.425 3.295 ;
        RECT  14.895 1.825 15.195 2.055 ;
        RECT  14.450 3.065 15.195 3.295 ;
        RECT  14.665 1.595 14.895 2.055 ;
        RECT  14.360 1.595 14.665 1.825 ;
        RECT  14.110 3.065 14.450 3.940 ;
        RECT  14.360 0.970 14.420 1.310 ;
        RECT  14.080 0.970 14.360 1.825 ;
        RECT  14.295 2.140 14.350 2.480 ;
        RECT  14.010 2.140 14.295 2.505 ;
        RECT  13.510 1.595 14.080 1.825 ;
        RECT  12.885 2.275 14.010 2.505 ;
        RECT  13.225 1.595 13.510 2.045 ;
        RECT  13.170 1.705 13.225 2.045 ;
        RECT  12.885 4.000 13.000 4.340 ;
        RECT  12.875 2.275 12.885 4.340 ;
        RECT  12.655 1.285 12.875 4.340 ;
        RECT  12.645 1.285 12.655 4.285 ;
        RECT  12.250 1.285 12.645 1.515 ;
        RECT  11.910 1.230 12.250 1.570 ;
        RECT  12.120 2.500 12.230 2.840 ;
        RECT  11.890 2.500 12.120 3.840 ;
        RECT  10.495 3.610 11.890 3.840 ;
        RECT  11.505 1.830 11.885 2.170 ;
        RECT  11.275 0.675 11.505 3.375 ;
        RECT  9.575 0.675 11.275 0.905 ;
        RECT  10.740 3.145 11.275 3.375 ;
        RECT  10.975 2.020 11.030 2.410 ;
        RECT  10.690 2.020 10.975 2.415 ;
        RECT  9.615 2.180 10.690 2.415 ;
        RECT  10.265 2.705 10.495 3.840 ;
        RECT  10.135 3.610 10.265 3.840 ;
        RECT  9.905 3.610 10.135 4.365 ;
        RECT  7.760 4.135 9.905 4.365 ;
        RECT  9.385 1.825 9.615 3.385 ;
        RECT  9.235 0.635 9.575 0.975 ;
        RECT  8.485 1.825 9.385 2.055 ;
        RECT  9.080 3.155 9.385 3.385 ;
        RECT  8.850 3.155 9.080 3.820 ;
        RECT  8.730 2.440 9.070 2.780 ;
        RECT  8.740 3.480 8.850 3.820 ;
        RECT  8.325 2.495 8.730 2.725 ;
        RECT  8.255 1.115 8.485 2.055 ;
        RECT  8.325 3.480 8.380 3.820 ;
        RECT  8.095 2.435 8.325 3.820 ;
        RECT  8.075 1.115 8.255 1.885 ;
        RECT  7.890 2.435 8.095 2.665 ;
        RECT  8.040 3.480 8.095 3.820 ;
        RECT  6.540 1.655 8.075 1.885 ;
        RECT  7.525 2.120 7.890 2.665 ;
        RECT  7.535 0.770 7.830 1.110 ;
        RECT  7.530 3.945 7.760 4.365 ;
        RECT  7.305 0.770 7.535 1.420 ;
        RECT  6.645 3.945 7.530 4.175 ;
        RECT  5.500 1.190 7.305 1.420 ;
        RECT  6.435 2.935 6.645 4.355 ;
        RECT  6.200 1.655 6.540 2.080 ;
        RECT  6.415 2.395 6.435 4.355 ;
        RECT  6.205 2.395 6.415 3.165 ;
        RECT  4.275 4.125 6.415 4.355 ;
        RECT  5.875 2.395 6.205 2.625 ;
        RECT  5.745 3.480 6.080 3.840 ;
        RECT  5.645 2.055 5.875 2.625 ;
        RECT  5.515 2.965 5.745 3.840 ;
        RECT  5.335 2.055 5.645 2.285 ;
        RECT  5.340 2.965 5.515 3.195 ;
        RECT  5.160 1.160 5.500 1.500 ;
        RECT  5.110 2.590 5.340 3.195 ;
        RECT  5.105 1.940 5.335 2.285 ;
        RECT  4.910 3.435 5.250 3.800 ;
        RECT  5.020 1.270 5.160 1.500 ;
        RECT  4.810 2.590 5.110 2.820 ;
        RECT  4.810 1.270 5.020 1.655 ;
        RECT  4.795 3.435 4.910 3.665 ;
        RECT  4.790 1.270 4.810 2.820 ;
        RECT  4.565 3.100 4.795 3.665 ;
        RECT  4.580 1.425 4.790 2.820 ;
        RECT  2.730 3.100 4.565 3.330 ;
        RECT  4.445 0.965 4.560 1.195 ;
        RECT  4.215 0.865 4.445 1.195 ;
        RECT  4.045 3.620 4.275 4.355 ;
        RECT  2.155 0.865 4.215 1.095 ;
        RECT  3.120 3.620 4.045 3.850 ;
        RECT  2.430 1.335 3.510 1.565 ;
        RECT  2.890 3.620 3.120 3.975 ;
        RECT  0.550 3.745 2.890 3.975 ;
        RECT  2.390 3.045 2.730 3.385 ;
        RECT  2.375 2.460 2.525 2.800 ;
        RECT  2.375 1.335 2.430 1.750 ;
        RECT  2.145 1.335 2.375 2.800 ;
        RECT  1.925 0.665 2.155 1.095 ;
        RECT  2.090 1.385 2.145 1.750 ;
        RECT  1.990 2.570 2.145 2.800 ;
        RECT  1.760 2.570 1.990 3.240 ;
        RECT  1.500 0.665 1.925 0.895 ;
        RECT  1.650 2.900 1.760 3.240 ;
        RECT  0.395 3.520 0.550 3.975 ;
        RECT  0.395 1.345 0.535 1.685 ;
        RECT  0.195 1.345 0.395 3.975 ;
        RECT  0.165 1.400 0.195 3.975 ;
    END
END SDFFRX1

MACRO SDFFNSRXL
    CLASS CORE ;
    FOREIGN SDFFNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.250 4.075 14.305 4.365 ;
        RECT  13.910 4.020 14.250 4.365 ;
        RECT  11.435 4.135 13.910 4.365 ;
        RECT  11.010 4.125 11.435 4.365 ;
        RECT  8.375 4.125 11.010 4.355 ;
        RECT  8.145 4.005 8.375 4.355 ;
        RECT  7.160 4.005 8.145 4.235 ;
        RECT  6.820 4.005 7.160 4.365 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 2.200 3.205 3.195 ;
        RECT  2.855 2.965 2.975 3.195 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.235 0.670 1.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.765 1.790 8.820 2.175 ;
        RECT  8.135 1.785 8.765 2.175 ;
        RECT  8.060 1.795 8.135 2.175 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.595 2.965 17.605 3.400 ;
        RECT  17.365 1.095 17.595 3.400 ;
        RECT  17.180 1.095 17.365 1.435 ;
        RECT  17.235 2.965 17.365 3.400 ;
        RECT  17.180 3.170 17.235 3.400 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.925 1.095 18.960 1.435 ;
        RECT  18.925 3.130 18.960 3.580 ;
        RECT  18.695 1.095 18.925 3.580 ;
        RECT  18.620 1.095 18.695 1.435 ;
        RECT  18.620 3.130 18.695 3.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.380 2.500 2.730 ;
        RECT  2.240 2.335 2.425 2.730 ;
        RECT  1.900 2.280 2.240 2.730 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  3.890 2.280 4.120 2.850 ;
        RECT  3.515 2.280 3.890 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.240 -0.400 19.140 0.400 ;
        RECT  17.900 -0.400 18.240 1.435 ;
        RECT  16.770 -0.400 17.900 0.400 ;
        RECT  16.430 -0.400 16.770 0.575 ;
        RECT  13.560 -0.400 16.430 0.400 ;
        RECT  13.220 -0.400 13.560 0.575 ;
        RECT  11.110 -0.400 13.220 0.400 ;
        RECT  10.770 -0.400 11.110 1.430 ;
        RECT  9.330 -0.400 10.770 0.400 ;
        RECT  8.990 -0.400 9.330 0.900 ;
        RECT  6.470 -0.400 8.990 0.400 ;
        RECT  6.130 -0.400 6.470 0.900 ;
        RECT  3.710 -0.400 6.130 0.400 ;
        RECT  3.370 -0.400 3.710 0.575 ;
        RECT  1.180 -0.400 3.370 0.400 ;
        RECT  0.840 -0.400 1.180 0.920 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.180 4.640 19.140 5.440 ;
        RECT  17.840 4.465 18.180 5.440 ;
        RECT  16.090 4.640 17.840 5.440 ;
        RECT  15.750 3.395 16.090 5.440 ;
        RECT  14.925 4.640 15.750 5.440 ;
        RECT  14.695 3.395 14.925 5.440 ;
        RECT  14.010 3.395 14.695 3.625 ;
        RECT  7.915 4.640 14.695 5.440 ;
        RECT  13.670 3.255 14.010 3.625 ;
        RECT  13.425 3.395 13.670 3.625 ;
        RECT  13.195 3.395 13.425 3.845 ;
        RECT  11.485 3.615 13.195 3.845 ;
        RECT  11.255 3.515 11.485 3.845 ;
        RECT  10.975 3.515 11.255 3.745 ;
        RECT  7.575 4.465 7.915 5.440 ;
        RECT  6.590 4.640 7.575 5.440 ;
        RECT  6.250 4.465 6.590 5.440 ;
        RECT  3.480 4.640 6.250 5.440 ;
        RECT  3.140 4.465 3.480 5.440 ;
        RECT  0.890 4.640 3.140 5.440 ;
        RECT  0.550 4.465 0.890 5.440 ;
        RECT  0.000 4.640 0.550 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.225 2.090 18.430 2.430 ;
        RECT  17.995 2.090 18.225 3.860 ;
        RECT  16.810 3.630 17.995 3.860 ;
        RECT  16.770 3.395 16.810 3.860 ;
        RECT  16.540 1.170 16.770 3.860 ;
        RECT  16.430 1.170 16.540 1.510 ;
        RECT  16.470 3.395 16.540 3.860 ;
        RECT  16.045 1.825 16.275 3.165 ;
        RECT  15.400 1.825 16.045 2.055 ;
        RECT  14.530 2.935 16.045 3.165 ;
        RECT  15.860 1.075 15.970 1.415 ;
        RECT  15.630 0.630 15.860 1.415 ;
        RECT  14.365 0.630 15.630 0.860 ;
        RECT  15.170 1.130 15.400 2.055 ;
        RECT  14.825 1.130 15.170 1.360 ;
        RECT  14.710 1.855 14.940 2.230 ;
        RECT  12.725 1.855 14.710 2.085 ;
        RECT  14.300 2.615 14.530 3.165 ;
        RECT  14.135 0.630 14.365 1.415 ;
        RECT  13.815 2.615 14.300 2.845 ;
        RECT  14.025 1.075 14.135 1.415 ;
        RECT  13.475 2.560 13.815 2.900 ;
        RECT  11.570 0.635 12.760 0.865 ;
        RECT  12.495 1.200 12.725 3.360 ;
        RECT  12.050 1.200 12.495 1.430 ;
        RECT  12.295 3.130 12.495 3.360 ;
        RECT  12.065 2.455 12.265 2.795 ;
        RECT  11.835 1.660 12.065 3.280 ;
        RECT  11.570 1.660 11.835 1.890 ;
        RECT  10.540 3.050 11.835 3.280 ;
        RECT  11.340 0.635 11.570 1.890 ;
        RECT  11.450 2.455 11.560 2.795 ;
        RECT  11.220 2.125 11.450 2.795 ;
        RECT  10.255 1.660 11.340 1.890 ;
        RECT  9.795 2.125 11.220 2.355 ;
        RECT  10.045 2.590 10.830 2.820 ;
        RECT  10.310 3.050 10.540 3.800 ;
        RECT  10.025 0.670 10.255 1.890 ;
        RECT  9.815 2.590 10.045 3.840 ;
        RECT  9.820 0.670 10.025 0.900 ;
        RECT  8.835 3.610 9.815 3.840 ;
        RECT  9.565 1.135 9.795 2.355 ;
        RECT  7.870 1.135 9.565 1.365 ;
        RECT  9.525 2.615 9.540 2.845 ;
        RECT  9.335 2.615 9.525 3.375 ;
        RECT  9.105 1.635 9.335 3.375 ;
        RECT  9.065 2.905 9.105 3.375 ;
        RECT  8.335 2.905 9.065 3.135 ;
        RECT  8.605 3.535 8.835 3.840 ;
        RECT  5.965 3.535 8.605 3.765 ;
        RECT  8.105 2.540 8.335 3.135 ;
        RECT  7.825 1.135 7.870 1.560 ;
        RECT  7.595 1.135 7.825 3.135 ;
        RECT  7.530 1.135 7.595 1.560 ;
        RECT  7.370 2.905 7.595 3.135 ;
        RECT  6.020 2.905 7.370 3.260 ;
        RECT  7.135 1.840 7.365 2.205 ;
        RECT  5.865 1.975 7.135 2.205 ;
        RECT  5.735 3.535 5.965 4.280 ;
        RECT  5.635 0.955 5.865 2.655 ;
        RECT  4.840 4.050 5.735 4.280 ;
        RECT  5.310 0.955 5.635 1.240 ;
        RECT  5.335 2.425 5.635 2.655 ;
        RECT  5.175 1.770 5.405 2.195 ;
        RECT  5.105 2.425 5.335 3.820 ;
        RECT  4.970 0.900 5.310 1.240 ;
        RECT  4.710 1.965 5.175 2.195 ;
        RECT  4.710 3.280 4.840 4.280 ;
        RECT  4.610 1.485 4.710 4.280 ;
        RECT  4.510 1.485 4.610 3.620 ;
        RECT  4.480 1.430 4.510 3.620 ;
        RECT  4.165 0.690 4.505 1.095 ;
        RECT  4.170 1.430 4.480 1.770 ;
        RECT  3.835 3.145 4.480 3.485 ;
        RECT  4.020 3.945 4.360 4.320 ;
        RECT  2.860 0.865 4.165 1.095 ;
        RECT  3.255 3.945 4.020 4.175 ;
        RECT  3.025 3.615 3.255 4.175 ;
        RECT  2.295 3.615 3.025 3.845 ;
        RECT  2.630 0.865 2.860 1.585 ;
        RECT  2.490 1.355 2.630 1.585 ;
        RECT  1.455 4.145 2.535 4.375 ;
        RECT  2.260 1.355 2.490 1.960 ;
        RECT  2.065 3.300 2.295 3.845 ;
        RECT  1.955 3.300 2.065 3.640 ;
        RECT  1.850 0.675 1.990 0.905 ;
        RECT  1.620 0.675 1.850 1.625 ;
        RECT  1.570 1.395 1.620 1.625 ;
        RECT  1.340 1.395 1.570 2.555 ;
        RECT  1.225 3.945 1.455 4.375 ;
        RECT  1.335 2.255 1.340 2.555 ;
        RECT  0.995 2.255 1.335 2.610 ;
        RECT  0.455 3.945 1.225 4.175 ;
        RECT  0.455 2.255 0.995 2.485 ;
        RECT  0.225 2.255 0.455 4.175 ;
    END
END SDFFNSRXL

MACRO SDFFNSRX4
    CLASS CORE ;
    FOREIGN SDFFNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSRXL ;
    SIZE 25.080 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.940 4.000 16.280 4.355 ;
        RECT  11.370 4.000 15.940 4.230 ;
        RECT  11.140 4.000 11.370 4.290 ;
        RECT  11.005 4.060 11.140 4.290 ;
        RECT  10.775 4.060 11.005 4.335 ;
        RECT  7.300 4.105 10.775 4.335 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.180 3.140 2.520 ;
        RECT  2.855 2.180 3.085 3.195 ;
        RECT  2.800 2.180 2.855 2.520 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 2.405 1.205 2.835 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.235 2.295 9.705 2.790 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.960 1.420 22.980 1.845 ;
        RECT  22.960 2.635 22.980 3.195 ;
        RECT  22.640 1.420 22.960 3.220 ;
        RECT  22.580 1.820 22.640 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.260 1.820 24.280 3.220 ;
        RECT  23.920 1.420 24.260 3.220 ;
        RECT  23.900 1.820 23.920 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 2.405 2.425 2.815 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 2.035 4.060 2.405 ;
        RECT  3.515 1.845 3.745 2.405 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.900 -0.400 25.080 0.400 ;
        RECT  24.560 -0.400 24.900 1.030 ;
        RECT  23.620 -0.400 24.560 0.400 ;
        RECT  23.280 -0.400 23.620 1.045 ;
        RECT  22.340 -0.400 23.280 0.400 ;
        RECT  22.000 -0.400 22.340 1.030 ;
        RECT  17.215 -0.400 22.000 0.400 ;
        RECT  16.875 -0.400 17.215 1.050 ;
        RECT  14.335 -0.400 16.875 0.400 ;
        RECT  13.995 -0.400 14.335 0.970 ;
        RECT  11.640 -0.400 13.995 0.400 ;
        RECT  11.410 -0.400 11.640 0.870 ;
        RECT  9.280 -0.400 11.410 0.400 ;
        RECT  8.940 -0.400 9.280 0.885 ;
        RECT  6.620 -0.400 8.940 0.400 ;
        RECT  6.280 -0.400 6.620 0.845 ;
        RECT  3.600 -0.400 6.280 0.400 ;
        RECT  3.260 -0.400 3.600 0.575 ;
        RECT  1.120 -0.400 3.260 0.400 ;
        RECT  0.780 -0.400 1.120 0.900 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.900 4.640 25.080 5.440 ;
        RECT  24.560 4.035 24.900 5.440 ;
        RECT  23.620 4.640 24.560 5.440 ;
        RECT  23.280 4.035 23.620 5.440 ;
        RECT  22.340 4.640 23.280 5.440 ;
        RECT  22.000 4.035 22.340 5.440 ;
        RECT  19.590 4.640 22.000 5.440 ;
        RECT  19.250 3.640 19.590 5.440 ;
        RECT  17.530 4.640 19.250 5.440 ;
        RECT  17.530 2.920 17.585 3.260 ;
        RECT  17.300 2.920 17.530 5.440 ;
        RECT  17.245 2.920 17.300 3.260 ;
        RECT  15.710 4.640 17.300 5.440 ;
        RECT  15.370 4.465 15.710 5.440 ;
        RECT  14.830 4.640 15.370 5.440 ;
        RECT  14.490 4.465 14.830 5.440 ;
        RECT  12.165 4.640 14.490 5.440 ;
        RECT  11.825 4.465 12.165 5.440 ;
        RECT  7.050 4.640 11.825 5.440 ;
        RECT  6.710 4.465 7.050 5.440 ;
        RECT  3.525 4.640 6.710 5.440 ;
        RECT  3.185 4.465 3.525 5.440 ;
        RECT  1.140 4.640 3.185 5.440 ;
        RECT  0.800 4.465 1.140 5.440 ;
        RECT  0.000 4.640 0.800 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  24.585 2.210 24.815 3.740 ;
        RECT  22.275 3.510 24.585 3.740 ;
        RECT  22.045 1.670 22.275 3.740 ;
        RECT  21.525 1.670 22.045 1.900 ;
        RECT  21.240 3.400 22.045 3.740 ;
        RECT  21.050 2.160 21.730 2.530 ;
        RECT  21.295 1.440 21.525 1.900 ;
        RECT  20.880 1.375 21.050 2.530 ;
        RECT  20.820 1.375 20.880 3.610 ;
        RECT  20.490 0.675 20.830 0.975 ;
        RECT  20.110 1.375 20.820 1.605 ;
        RECT  20.650 2.300 20.820 3.610 ;
        RECT  20.540 3.085 20.650 3.610 ;
        RECT  20.420 1.835 20.590 2.065 ;
        RECT  18.310 3.085 20.540 3.315 ;
        RECT  19.390 0.675 20.490 0.905 ;
        RECT  20.190 1.835 20.420 2.155 ;
        RECT  18.440 1.925 20.190 2.155 ;
        RECT  19.740 1.185 20.110 1.605 ;
        RECT  18.765 1.375 19.740 1.605 ;
        RECT  19.050 0.675 19.390 1.050 ;
        RECT  17.940 0.675 19.050 0.905 ;
        RECT  18.535 1.140 18.765 1.605 ;
        RECT  18.325 1.140 18.535 1.370 ;
        RECT  18.085 1.895 18.440 2.155 ;
        RECT  18.200 3.085 18.310 3.600 ;
        RECT  17.970 2.455 18.200 3.600 ;
        RECT  15.860 1.925 18.085 2.155 ;
        RECT  16.865 2.455 17.970 2.685 ;
        RECT  17.830 0.675 17.940 1.290 ;
        RECT  17.710 0.675 17.830 1.605 ;
        RECT  17.600 0.950 17.710 1.605 ;
        RECT  16.495 1.375 17.600 1.605 ;
        RECT  16.840 3.535 17.070 4.410 ;
        RECT  16.635 2.455 16.865 3.305 ;
        RECT  10.835 3.535 16.840 3.765 ;
        RECT  16.525 2.810 16.635 3.305 ;
        RECT  14.500 3.075 16.525 3.305 ;
        RECT  16.265 0.970 16.495 1.605 ;
        RECT  16.155 0.970 16.265 1.310 ;
        RECT  15.655 0.865 15.860 2.155 ;
        RECT  15.630 0.865 15.655 2.845 ;
        RECT  15.355 0.865 15.630 1.095 ;
        RECT  15.425 1.925 15.630 2.845 ;
        RECT  13.695 1.925 15.425 2.155 ;
        RECT  15.060 1.350 15.400 1.690 ;
        RECT  14.500 2.385 15.160 2.615 ;
        RECT  13.535 1.350 15.060 1.580 ;
        RECT  14.270 2.385 14.500 3.305 ;
        RECT  13.465 1.815 13.695 3.135 ;
        RECT  13.305 0.675 13.535 1.580 ;
        RECT  13.015 1.815 13.465 2.045 ;
        RECT  13.155 2.905 13.465 3.135 ;
        RECT  12.380 0.675 13.305 0.905 ;
        RECT  12.380 2.275 13.230 2.505 ;
        RECT  12.785 1.220 13.015 2.045 ;
        RECT  12.675 1.220 12.785 1.560 ;
        RECT  12.150 0.675 12.380 3.195 ;
        RECT  11.295 2.965 12.150 3.195 ;
        RECT  11.690 1.530 11.920 2.170 ;
        RECT  11.180 1.530 11.690 1.760 ;
        RECT  11.065 2.275 11.295 3.195 ;
        RECT  10.950 0.840 11.180 1.760 ;
        RECT  10.720 2.275 11.065 2.505 ;
        RECT  9.970 0.840 10.950 1.070 ;
        RECT  10.605 3.085 10.835 3.765 ;
        RECT  10.490 1.300 10.720 2.505 ;
        RECT  10.220 3.085 10.605 3.315 ;
        RECT  10.450 2.145 10.490 2.505 ;
        RECT  10.320 3.605 10.375 3.835 ;
        RECT  10.090 3.605 10.320 3.840 ;
        RECT  9.990 1.625 10.220 3.315 ;
        RECT  6.275 3.610 10.090 3.840 ;
        RECT  9.620 1.625 9.990 1.855 ;
        RECT  8.810 3.085 9.990 3.315 ;
        RECT  9.740 0.840 9.970 1.395 ;
        RECT  8.030 1.165 9.740 1.395 ;
        RECT  8.580 2.280 8.810 3.315 ;
        RECT  8.470 2.280 8.580 2.620 ;
        RECT  7.800 1.165 8.030 3.375 ;
        RECT  7.660 1.165 7.800 1.505 ;
        RECT  6.655 3.145 7.800 3.375 ;
        RECT  7.230 1.900 7.570 2.240 ;
        RECT  5.960 1.955 7.230 2.185 ;
        RECT  6.315 3.035 6.655 3.375 ;
        RECT  6.045 3.610 6.275 4.410 ;
        RECT  5.230 4.180 6.045 4.410 ;
        RECT  5.730 0.745 5.960 3.080 ;
        RECT  5.620 0.745 5.730 1.030 ;
        RECT  5.690 2.850 5.730 3.080 ;
        RECT  5.460 2.850 5.690 3.920 ;
        RECT  5.280 0.690 5.620 1.030 ;
        RECT  4.615 1.940 5.500 2.280 ;
        RECT  5.000 3.045 5.230 4.410 ;
        RECT  4.890 3.045 5.000 3.385 ;
        RECT  4.560 0.730 4.900 1.070 ;
        RECT  4.615 3.045 4.890 3.360 ;
        RECT  4.540 3.735 4.770 4.120 ;
        RECT  4.385 1.490 4.615 3.360 ;
        RECT  2.605 0.805 4.560 1.035 ;
        RECT  3.585 3.735 4.540 3.965 ;
        RECT  4.060 1.490 4.385 1.720 ;
        RECT  3.945 3.020 4.385 3.360 ;
        RECT  3.355 3.605 3.585 3.965 ;
        RECT  2.400 3.605 3.355 3.835 ;
        RECT  1.685 4.125 2.750 4.355 ;
        RECT  2.375 0.805 2.605 1.590 ;
        RECT  2.170 3.130 2.400 3.835 ;
        RECT  2.100 1.250 2.375 1.590 ;
        RECT  2.060 3.130 2.170 3.470 ;
        RECT  1.455 3.185 1.685 4.355 ;
        RECT  0.520 1.865 1.470 2.095 ;
        RECT  0.520 3.185 1.455 3.415 ;
        RECT  0.405 1.390 0.520 2.095 ;
        RECT  0.405 3.130 0.520 3.470 ;
        RECT  0.180 1.390 0.405 3.470 ;
        RECT  0.175 1.400 0.180 3.470 ;
    END
END SDFFNSRX4

MACRO SDFFNSRX2
    CLASS CORE ;
    FOREIGN SDFFNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.250 4.070 14.305 4.365 ;
        RECT  13.910 4.015 14.250 4.365 ;
        RECT  8.375 4.135 13.910 4.365 ;
        RECT  8.145 4.005 8.375 4.365 ;
        RECT  7.340 4.005 8.145 4.235 ;
        RECT  7.110 4.005 7.340 4.365 ;
        RECT  7.045 4.085 7.110 4.365 ;
        RECT  6.820 4.135 7.045 4.365 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.230 2.200 3.265 2.540 ;
        RECT  3.000 2.200 3.230 3.195 ;
        RECT  2.925 2.200 3.000 2.540 ;
        RECT  2.855 2.965 3.000 3.195 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.690 2.820 1.180 3.340 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.425 1.785 9.100 2.175 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.680 1.440 17.855 2.970 ;
        RECT  17.625 1.440 17.680 3.080 ;
        RECT  17.340 1.440 17.625 1.780 ;
        RECT  17.375 2.740 17.625 3.195 ;
        RECT  17.340 2.740 17.375 3.080 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.765 1.440 18.995 3.195 ;
        RECT  18.620 1.440 18.765 1.780 ;
        RECT  18.695 2.740 18.765 3.195 ;
        RECT  18.620 2.740 18.695 3.080 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 2.280 2.500 2.730 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  4.230 2.270 4.480 2.660 ;
        RECT  3.890 2.270 4.230 2.715 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.320 -0.400 19.140 0.400 ;
        RECT  17.980 -0.400 18.320 1.030 ;
        RECT  16.835 -0.400 17.980 0.400 ;
        RECT  16.495 -0.400 16.835 0.575 ;
        RECT  13.835 -0.400 16.495 0.400 ;
        RECT  13.495 -0.400 13.835 0.575 ;
        RECT  11.335 -0.400 13.495 0.400 ;
        RECT  10.995 -0.400 11.335 1.370 ;
        RECT  9.575 -0.400 10.995 0.400 ;
        RECT  9.235 -0.400 9.575 0.900 ;
        RECT  6.475 -0.400 9.235 0.400 ;
        RECT  6.135 -0.400 6.475 0.900 ;
        RECT  3.710 -0.400 6.135 0.400 ;
        RECT  3.370 -0.400 3.710 0.575 ;
        RECT  1.155 -0.400 3.370 0.400 ;
        RECT  0.815 -0.400 1.155 0.970 ;
        RECT  0.000 -0.400 0.815 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.320 4.640 19.140 5.440 ;
        RECT  17.980 4.090 18.320 5.440 ;
        RECT  16.010 4.640 17.980 5.440 ;
        RECT  15.670 3.560 16.010 5.440 ;
        RECT  14.925 4.640 15.670 5.440 ;
        RECT  14.695 3.485 14.925 5.440 ;
        RECT  13.425 3.485 14.695 3.715 ;
        RECT  7.915 4.640 14.695 5.440 ;
        RECT  13.195 3.485 13.425 3.845 ;
        RECT  11.485 3.615 13.195 3.845 ;
        RECT  11.255 3.515 11.485 3.845 ;
        RECT  11.015 3.515 11.255 3.745 ;
        RECT  7.575 4.465 7.915 5.440 ;
        RECT  6.590 4.640 7.575 5.440 ;
        RECT  6.250 4.465 6.590 5.440 ;
        RECT  3.480 4.640 6.250 5.440 ;
        RECT  3.140 4.465 3.480 5.440 ;
        RECT  0.890 4.640 3.140 5.440 ;
        RECT  0.550 4.465 0.890 5.440 ;
        RECT  0.000 4.640 0.550 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.315 2.090 18.535 2.430 ;
        RECT  18.085 2.090 18.315 3.830 ;
        RECT  17.070 3.600 18.085 3.830 ;
        RECT  16.845 1.225 17.070 3.830 ;
        RECT  16.840 1.170 16.845 3.830 ;
        RECT  16.505 1.170 16.840 1.510 ;
        RECT  16.735 3.600 16.840 3.830 ;
        RECT  16.395 3.600 16.735 4.005 ;
        RECT  16.380 2.300 16.490 2.640 ;
        RECT  16.150 1.825 16.380 3.165 ;
        RECT  15.385 1.825 16.150 2.055 ;
        RECT  14.335 2.935 16.150 3.165 ;
        RECT  15.695 0.760 16.035 1.120 ;
        RECT  14.595 0.760 15.695 0.990 ;
        RECT  15.155 1.220 15.385 2.055 ;
        RECT  14.975 1.220 15.155 1.560 ;
        RECT  14.580 1.890 14.920 2.230 ;
        RECT  14.255 0.760 14.595 1.120 ;
        RECT  13.585 1.890 14.580 2.120 ;
        RECT  14.105 2.670 14.335 3.165 ;
        RECT  13.590 2.670 14.105 2.900 ;
        RECT  13.250 2.560 13.590 2.900 ;
        RECT  13.355 1.335 13.585 2.120 ;
        RECT  12.935 1.335 13.355 1.565 ;
        RECT  12.045 0.735 13.065 0.965 ;
        RECT  12.705 1.335 12.935 3.325 ;
        RECT  12.615 1.335 12.705 1.620 ;
        RECT  12.295 3.095 12.705 3.325 ;
        RECT  12.275 1.280 12.615 1.620 ;
        RECT  12.045 2.470 12.370 2.810 ;
        RECT  11.815 0.735 12.045 3.285 ;
        RECT  10.480 1.600 11.815 1.830 ;
        RECT  10.635 3.055 11.815 3.285 ;
        RECT  11.310 2.060 11.540 2.515 ;
        RECT  10.020 2.060 11.310 2.290 ;
        RECT  10.060 2.525 10.755 2.755 ;
        RECT  10.405 3.055 10.635 3.800 ;
        RECT  10.250 0.630 10.480 1.830 ;
        RECT  10.295 3.460 10.405 3.800 ;
        RECT  10.045 0.630 10.250 0.860 ;
        RECT  9.830 2.525 10.060 3.890 ;
        RECT  9.790 1.135 10.020 2.290 ;
        RECT  8.835 3.660 9.830 3.890 ;
        RECT  7.950 1.135 9.790 1.365 ;
        RECT  9.330 1.600 9.560 3.375 ;
        RECT  9.220 2.480 9.330 3.375 ;
        RECT  9.065 2.905 9.220 3.375 ;
        RECT  8.380 2.905 9.065 3.135 ;
        RECT  8.605 3.520 8.835 3.890 ;
        RECT  5.930 3.520 8.605 3.750 ;
        RECT  8.150 2.540 8.380 3.135 ;
        RECT  7.920 1.120 7.950 1.460 ;
        RECT  7.690 1.120 7.920 3.135 ;
        RECT  7.610 1.120 7.690 1.460 ;
        RECT  7.370 2.905 7.690 3.135 ;
        RECT  7.215 1.840 7.445 2.205 ;
        RECT  6.325 2.905 7.370 3.260 ;
        RECT  5.865 1.975 7.215 2.205 ;
        RECT  6.095 2.510 6.325 3.260 ;
        RECT  5.700 3.520 5.930 4.325 ;
        RECT  5.635 0.955 5.865 2.965 ;
        RECT  4.785 4.095 5.700 4.325 ;
        RECT  5.310 0.955 5.635 1.240 ;
        RECT  5.470 2.735 5.635 2.965 ;
        RECT  5.240 2.735 5.470 3.820 ;
        RECT  4.945 1.770 5.405 2.115 ;
        RECT  4.970 0.900 5.310 1.240 ;
        RECT  5.105 3.480 5.240 3.820 ;
        RECT  4.790 1.510 4.945 3.125 ;
        RECT  4.785 1.510 4.790 3.535 ;
        RECT  4.715 1.510 4.785 4.325 ;
        RECT  4.510 1.510 4.715 1.740 ;
        RECT  4.560 2.895 4.715 4.325 ;
        RECT  4.555 3.250 4.560 4.325 ;
        RECT  4.495 3.250 4.555 3.645 ;
        RECT  4.170 1.400 4.510 1.740 ;
        RECT  4.290 0.685 4.505 0.915 ;
        RECT  3.835 3.250 4.495 3.590 ;
        RECT  4.075 3.945 4.305 4.320 ;
        RECT  4.060 0.685 4.290 1.095 ;
        RECT  3.255 3.945 4.075 4.175 ;
        RECT  2.860 0.865 4.060 1.095 ;
        RECT  3.025 3.615 3.255 4.175 ;
        RECT  2.295 3.615 3.025 3.845 ;
        RECT  2.630 0.865 2.860 1.585 ;
        RECT  2.490 1.355 2.630 1.585 ;
        RECT  1.455 4.145 2.535 4.375 ;
        RECT  2.260 1.355 2.490 1.960 ;
        RECT  2.065 3.300 2.295 3.845 ;
        RECT  1.955 3.300 2.065 3.640 ;
        RECT  1.840 0.685 1.985 0.915 ;
        RECT  1.610 0.685 1.840 1.625 ;
        RECT  1.570 1.395 1.610 1.625 ;
        RECT  1.340 1.395 1.570 2.500 ;
        RECT  1.225 3.945 1.455 4.375 ;
        RECT  1.230 2.160 1.340 2.500 ;
        RECT  0.455 2.270 1.230 2.500 ;
        RECT  0.455 3.945 1.225 4.175 ;
        RECT  0.225 2.270 0.455 4.175 ;
    END
END SDFFNSRX2

MACRO SDFFNSRX1
    CLASS CORE ;
    FOREIGN SDFFNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.720 3.980 14.015 4.320 ;
        RECT  13.675 3.980 13.720 4.365 ;
        RECT  13.415 4.035 13.675 4.365 ;
        RECT  11.435 4.135 13.415 4.365 ;
        RECT  11.010 4.125 11.435 4.365 ;
        RECT  8.140 4.125 11.010 4.355 ;
        RECT  7.910 4.005 8.140 4.355 ;
        RECT  6.925 4.005 7.910 4.235 ;
        RECT  6.585 4.005 6.925 4.345 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.730 2.605 3.210 3.220 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.820 0.880 3.340 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 1.785 8.830 2.175 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.595 2.965 17.605 3.400 ;
        RECT  17.365 1.095 17.595 3.400 ;
        RECT  17.180 1.095 17.365 1.435 ;
        RECT  17.050 3.170 17.365 3.400 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.730 1.050 18.960 3.780 ;
        RECT  18.620 1.050 18.730 1.390 ;
        RECT  18.695 2.955 18.730 3.780 ;
        RECT  18.620 3.125 18.695 3.780 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.860 2.280 2.500 2.730 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.380 4.000 2.970 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.240 -0.400 19.140 0.400 ;
        RECT  17.900 -0.400 18.240 1.390 ;
        RECT  16.800 -0.400 17.900 0.400 ;
        RECT  16.460 -0.400 16.800 0.575 ;
        RECT  13.760 -0.400 16.460 0.400 ;
        RECT  13.420 -0.400 13.760 0.575 ;
        RECT  11.175 -0.400 13.420 0.400 ;
        RECT  10.835 -0.400 11.175 1.380 ;
        RECT  9.215 -0.400 10.835 0.400 ;
        RECT  8.875 -0.400 9.215 0.900 ;
        RECT  6.490 -0.400 8.875 0.400 ;
        RECT  6.150 -0.400 6.490 0.900 ;
        RECT  3.730 -0.400 6.150 0.400 ;
        RECT  3.390 -0.400 3.730 0.575 ;
        RECT  1.145 -0.400 3.390 0.400 ;
        RECT  0.805 -0.400 1.145 1.000 ;
        RECT  0.000 -0.400 0.805 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.200 4.640 19.140 5.440 ;
        RECT  17.860 4.090 18.200 5.440 ;
        RECT  15.855 4.640 17.860 5.440 ;
        RECT  15.515 3.395 15.855 5.440 ;
        RECT  14.690 4.640 15.515 5.440 ;
        RECT  14.460 3.390 14.690 5.440 ;
        RECT  13.160 3.390 14.460 3.620 ;
        RECT  7.680 4.640 14.460 5.440 ;
        RECT  12.930 3.390 13.160 3.845 ;
        RECT  11.080 3.615 12.930 3.845 ;
        RECT  10.740 3.455 11.080 3.845 ;
        RECT  7.340 4.465 7.680 5.440 ;
        RECT  6.355 4.640 7.340 5.440 ;
        RECT  6.015 4.465 6.355 5.440 ;
        RECT  3.270 4.640 6.015 5.440 ;
        RECT  2.930 4.465 3.270 5.440 ;
        RECT  0.700 4.640 2.930 5.440 ;
        RECT  0.360 4.465 0.700 5.440 ;
        RECT  0.000 4.640 0.360 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.320 2.090 18.480 2.430 ;
        RECT  18.090 2.090 18.320 3.860 ;
        RECT  16.820 3.630 18.090 3.860 ;
        RECT  16.590 1.170 16.820 3.860 ;
        RECT  16.480 1.170 16.590 1.510 ;
        RECT  16.235 3.395 16.590 3.735 ;
        RECT  16.225 2.300 16.335 2.640 ;
        RECT  15.995 1.825 16.225 3.160 ;
        RECT  15.890 1.055 16.000 1.395 ;
        RECT  15.305 1.825 15.995 2.055 ;
        RECT  14.100 2.930 15.995 3.160 ;
        RECT  15.660 0.630 15.890 1.395 ;
        RECT  14.560 0.630 15.660 0.860 ;
        RECT  15.075 1.090 15.305 2.055 ;
        RECT  14.940 1.090 15.075 1.320 ;
        RECT  14.460 1.890 14.800 2.230 ;
        RECT  14.330 0.630 14.560 1.395 ;
        RECT  13.350 1.890 14.460 2.120 ;
        RECT  14.220 1.055 14.330 1.395 ;
        RECT  13.870 2.670 14.100 3.160 ;
        RECT  13.420 2.670 13.870 2.900 ;
        RECT  13.080 2.560 13.420 2.900 ;
        RECT  13.120 1.175 13.350 2.120 ;
        RECT  12.700 1.175 13.120 1.405 ;
        RECT  11.825 0.715 12.985 0.945 ;
        RECT  12.470 1.175 12.700 3.360 ;
        RECT  12.115 1.175 12.470 1.405 ;
        RECT  12.060 3.130 12.470 3.360 ;
        RECT  11.845 2.485 12.155 2.825 ;
        RECT  11.825 1.615 11.845 2.825 ;
        RECT  11.595 0.715 11.825 3.225 ;
        RECT  10.320 1.615 11.595 1.845 ;
        RECT  10.305 2.995 11.595 3.225 ;
        RECT  11.130 2.075 11.360 2.605 ;
        RECT  9.860 2.075 11.130 2.305 ;
        RECT  9.825 2.535 10.655 2.765 ;
        RECT  10.090 0.675 10.320 1.845 ;
        RECT  10.075 2.995 10.305 3.740 ;
        RECT  9.880 0.675 10.090 0.905 ;
        RECT  9.630 1.135 9.860 2.305 ;
        RECT  9.595 2.535 9.825 3.845 ;
        RECT  7.890 1.135 9.630 1.365 ;
        RECT  8.600 3.615 9.595 3.845 ;
        RECT  9.345 1.635 9.400 1.975 ;
        RECT  9.115 1.635 9.345 3.375 ;
        RECT  9.060 1.635 9.115 1.975 ;
        RECT  9.005 2.480 9.115 3.375 ;
        RECT  8.830 2.905 9.005 3.375 ;
        RECT  8.190 2.905 8.830 3.135 ;
        RECT  8.370 3.515 8.600 3.845 ;
        RECT  5.720 3.515 8.370 3.745 ;
        RECT  7.960 2.540 8.190 3.135 ;
        RECT  7.730 1.120 7.890 1.460 ;
        RECT  7.500 1.120 7.730 3.135 ;
        RECT  7.135 2.905 7.500 3.135 ;
        RECT  7.040 2.180 7.270 2.535 ;
        RECT  5.900 2.905 7.135 3.260 ;
        RECT  5.920 2.180 7.040 2.410 ;
        RECT  5.690 0.955 5.920 2.650 ;
        RECT  5.490 3.515 5.720 4.320 ;
        RECT  5.330 0.955 5.690 1.240 ;
        RECT  5.155 2.420 5.690 2.650 ;
        RECT  4.585 4.090 5.490 4.320 ;
        RECT  5.230 1.770 5.460 2.185 ;
        RECT  4.990 0.900 5.330 1.240 ;
        RECT  4.530 1.955 5.230 2.185 ;
        RECT  4.925 2.420 5.155 3.820 ;
        RECT  4.815 3.480 4.925 3.820 ;
        RECT  4.475 3.250 4.585 4.320 ;
        RECT  4.190 0.630 4.530 1.095 ;
        RECT  4.475 1.400 4.530 2.185 ;
        RECT  4.355 1.400 4.475 4.320 ;
        RECT  4.245 1.400 4.355 3.645 ;
        RECT  4.190 1.400 4.245 1.740 ;
        RECT  3.690 3.250 4.245 3.590 ;
        RECT  2.625 0.865 4.190 1.095 ;
        RECT  3.785 3.945 4.125 4.380 ;
        RECT  3.020 3.945 3.785 4.175 ;
        RECT  2.790 3.615 3.020 4.175 ;
        RECT  2.060 3.615 2.790 3.845 ;
        RECT  2.395 0.865 2.625 1.740 ;
        RECT  2.230 1.400 2.395 1.740 ;
        RECT  1.340 4.145 2.300 4.375 ;
        RECT  1.830 3.295 2.060 3.845 ;
        RECT  1.770 0.715 2.010 0.945 ;
        RECT  1.720 3.295 1.830 3.635 ;
        RECT  1.540 0.715 1.770 1.460 ;
        RECT  1.340 1.230 1.540 1.460 ;
        RECT  1.340 2.190 1.455 2.530 ;
        RECT  1.110 1.230 1.340 4.375 ;
    END
END SDFFNSRX1

MACRO SDFFNSXL
    CLASS CORE ;
    FOREIGN SDFFNSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.575 3.475 13.190 3.915 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 2.150 3.810 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.700 1.860 2.250 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.965 0.865 14.985 3.755 ;
        RECT  14.755 0.865 14.965 4.010 ;
        RECT  14.340 0.865 14.755 1.095 ;
        RECT  14.735 3.525 14.755 4.010 ;
        RECT  14.380 3.780 14.735 4.010 ;
        RECT  14.340 3.780 14.380 4.085 ;
        RECT  14.000 0.715 14.340 1.095 ;
        RECT  14.000 3.780 14.340 4.195 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.625 1.250 15.660 1.845 ;
        RECT  15.625 3.095 15.660 3.435 ;
        RECT  15.395 1.250 15.625 3.435 ;
        RECT  15.320 1.250 15.395 1.820 ;
        RECT  15.320 3.095 15.395 3.435 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.345 4.405 2.075 ;
        RECT  4.100 1.345 4.175 1.820 ;
        RECT  4.015 1.345 4.100 1.685 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.280 1.180 2.700 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.100 -0.400 15.840 0.400 ;
        RECT  14.760 -0.400 15.100 0.575 ;
        RECT  13.560 -0.400 14.760 0.400 ;
        RECT  13.220 -0.400 13.560 0.575 ;
        RECT  11.680 -0.400 13.220 0.400 ;
        RECT  11.340 -0.400 11.680 0.575 ;
        RECT  9.110 -0.400 11.340 0.400 ;
        RECT  8.880 -0.400 9.110 1.135 ;
        RECT  6.800 -0.400 8.880 0.400 ;
        RECT  6.460 -0.400 6.800 1.065 ;
        RECT  3.275 -0.400 6.460 0.400 ;
        RECT  2.935 -0.400 3.275 0.575 ;
        RECT  1.200 -0.400 2.935 0.400 ;
        RECT  0.860 -0.400 1.200 0.575 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.100 4.640 15.840 5.440 ;
        RECT  14.760 4.465 15.100 5.440 ;
        RECT  13.580 4.640 14.760 5.440 ;
        RECT  13.240 4.465 13.580 5.440 ;
        RECT  12.320 4.640 13.240 5.440 ;
        RECT  11.980 4.140 12.320 5.440 ;
        RECT  9.800 4.640 11.980 5.440 ;
        RECT  9.460 3.755 9.800 5.440 ;
        RECT  8.340 4.640 9.460 5.440 ;
        RECT  8.000 4.160 8.340 5.440 ;
        RECT  7.045 4.640 8.000 5.440 ;
        RECT  6.705 4.465 7.045 5.440 ;
        RECT  3.660 4.640 6.705 5.440 ;
        RECT  3.320 4.155 3.660 5.440 ;
        RECT  1.080 4.640 3.320 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.295 1.430 14.525 3.190 ;
        RECT  14.020 1.430 14.295 1.770 ;
        RECT  14.000 2.960 14.295 3.190 ;
        RECT  13.570 2.140 13.910 2.480 ;
        RECT  13.155 2.195 13.570 2.425 ;
        RECT  12.925 1.620 13.155 3.245 ;
        RECT  12.380 1.620 12.925 1.850 ;
        RECT  12.660 2.905 12.925 3.245 ;
        RECT  11.195 2.290 12.670 2.520 ;
        RECT  12.040 1.190 12.380 1.850 ;
        RECT  11.850 1.620 12.040 1.850 ;
        RECT  11.510 1.620 11.850 1.960 ;
        RECT  10.965 1.300 11.195 3.890 ;
        RECT  10.520 1.300 10.965 1.530 ;
        RECT  10.740 3.550 10.965 3.890 ;
        RECT  9.855 0.645 10.930 0.875 ;
        RECT  9.855 2.550 10.735 2.890 ;
        RECT  10.180 1.190 10.520 1.530 ;
        RECT  9.625 0.645 9.855 2.890 ;
        RECT  8.650 1.370 9.625 1.600 ;
        RECT  9.100 2.660 9.625 2.890 ;
        RECT  9.055 1.830 9.395 2.170 ;
        RECT  8.870 2.660 9.100 3.470 ;
        RECT  8.435 1.885 9.055 2.115 ;
        RECT  8.760 3.130 8.870 3.470 ;
        RECT  8.585 3.700 8.815 4.040 ;
        RECT  8.420 0.695 8.650 1.600 ;
        RECT  6.250 3.700 8.585 3.930 ;
        RECT  8.205 1.885 8.435 3.415 ;
        RECT  7.295 0.630 8.420 0.925 ;
        RECT  8.190 1.885 8.205 2.115 ;
        RECT  7.105 3.185 8.205 3.415 ;
        RECT  7.960 1.450 8.190 2.115 ;
        RECT  7.625 2.400 7.965 2.740 ;
        RECT  7.395 1.295 7.625 2.630 ;
        RECT  5.435 1.295 7.395 1.525 ;
        RECT  6.875 2.090 7.105 3.415 ;
        RECT  6.735 2.090 6.875 2.320 ;
        RECT  6.395 1.980 6.735 2.320 ;
        RECT  6.020 2.570 6.250 4.055 ;
        RECT  5.945 2.570 6.020 2.800 ;
        RECT  5.300 3.825 6.020 4.055 ;
        RECT  5.715 1.755 5.945 2.800 ;
        RECT  5.480 3.180 5.780 3.520 ;
        RECT  5.460 1.755 5.715 1.985 ;
        RECT  5.250 2.595 5.480 3.520 ;
        RECT  5.145 0.815 5.435 1.525 ;
        RECT  4.960 3.825 5.300 4.170 ;
        RECT  5.145 2.595 5.250 2.825 ;
        RECT  5.095 0.815 5.145 2.825 ;
        RECT  4.915 1.295 5.095 2.825 ;
        RECT  4.680 3.110 5.020 3.450 ;
        RECT  4.145 3.825 4.960 4.055 ;
        RECT  2.540 3.170 4.680 3.400 ;
        RECT  4.295 0.740 4.635 1.080 ;
        RECT  1.900 0.850 4.295 1.080 ;
        RECT  3.915 3.690 4.145 4.055 ;
        RECT  2.970 3.690 3.915 3.920 ;
        RECT  3.260 1.345 3.600 1.685 ;
        RECT  2.430 1.440 3.260 1.670 ;
        RECT  2.740 3.690 2.970 4.175 ;
        RECT  2.375 2.490 2.780 2.830 ;
        RECT  0.520 3.945 2.740 4.175 ;
        RECT  2.200 3.060 2.540 3.400 ;
        RECT  2.375 1.440 2.430 1.780 ;
        RECT  2.145 1.440 2.375 2.830 ;
        RECT  2.090 1.440 2.145 1.780 ;
        RECT  1.840 2.600 2.145 2.830 ;
        RECT  1.560 0.640 1.900 1.080 ;
        RECT  1.610 2.600 1.840 3.610 ;
        RECT  1.500 3.270 1.610 3.610 ;
        RECT  0.395 1.195 0.540 1.535 ;
        RECT  0.395 3.270 0.520 4.175 ;
        RECT  0.290 1.195 0.395 4.175 ;
        RECT  0.165 1.195 0.290 3.610 ;
    END
END SDFFNSXL

MACRO SDFFNSX4
    CLASS CORE ;
    FOREIGN SDFFNSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.110 4.010 7.730 4.390 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.005 3.210 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.440 1.700 1.840 2.410 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.660 2.875 19.675 3.215 ;
        RECT  19.440 1.200 19.660 3.215 ;
        RECT  19.335 0.715 19.440 3.215 ;
        RECT  19.280 0.715 19.335 2.660 ;
        RECT  19.100 0.715 19.280 1.655 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.980 0.955 20.990 2.700 ;
        RECT  20.880 0.955 20.980 3.220 ;
        RECT  20.600 0.760 20.880 3.220 ;
        RECT  20.595 0.760 20.600 3.160 ;
        RECT  20.540 0.760 20.595 1.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.230 1.410 4.570 2.090 ;
        RECT  4.175 1.835 4.230 2.075 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 2.055 1.170 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.600 -0.400 21.780 0.400 ;
        RECT  21.260 -0.400 21.600 1.565 ;
        RECT  20.160 -0.400 21.260 0.400 ;
        RECT  19.820 -0.400 20.160 0.960 ;
        RECT  18.680 -0.400 19.820 0.400 ;
        RECT  18.340 -0.400 18.680 0.915 ;
        RECT  17.420 -0.400 18.340 0.400 ;
        RECT  17.080 -0.400 17.420 1.190 ;
        RECT  14.815 -0.400 17.080 0.400 ;
        RECT  14.475 -0.400 14.815 0.575 ;
        RECT  12.740 -0.400 14.475 0.400 ;
        RECT  12.400 -0.400 12.740 0.575 ;
        RECT  10.060 -0.400 12.400 0.400 ;
        RECT  9.720 -0.400 10.060 1.080 ;
        RECT  7.015 -0.400 9.720 0.400 ;
        RECT  6.675 -0.400 7.015 1.215 ;
        RECT  3.490 -0.400 6.675 0.400 ;
        RECT  3.150 -0.400 3.490 0.575 ;
        RECT  1.395 -0.400 3.150 0.400 ;
        RECT  1.055 -0.400 1.395 0.575 ;
        RECT  0.000 -0.400 1.055 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.595 4.640 21.780 5.440 ;
        RECT  21.255 4.055 21.595 5.440 ;
        RECT  20.315 4.640 21.255 5.440 ;
        RECT  19.975 4.015 20.315 5.440 ;
        RECT  19.035 4.640 19.975 5.440 ;
        RECT  18.695 4.055 19.035 5.440 ;
        RECT  17.610 4.640 18.695 5.440 ;
        RECT  17.270 3.520 17.610 5.440 ;
        RECT  16.170 4.640 17.270 5.440 ;
        RECT  15.830 3.520 16.170 5.440 ;
        RECT  14.690 4.640 15.830 5.440 ;
        RECT  14.350 3.960 14.690 5.440 ;
        RECT  12.620 4.640 14.350 5.440 ;
        RECT  12.280 3.380 12.620 5.440 ;
        RECT  10.020 4.640 12.280 5.440 ;
        RECT  9.680 3.330 10.020 5.440 ;
        RECT  8.360 4.640 9.680 5.440 ;
        RECT  8.020 4.195 8.360 5.440 ;
        RECT  6.870 4.640 8.020 5.440 ;
        RECT  6.530 4.150 6.870 5.440 ;
        RECT  3.665 4.640 6.530 5.440 ;
        RECT  3.325 4.195 3.665 5.440 ;
        RECT  1.080 4.640 3.325 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.285 2.060 21.515 3.725 ;
        RECT  18.755 3.495 21.285 3.725 ;
        RECT  18.525 1.620 18.755 3.725 ;
        RECT  18.140 1.620 18.525 1.850 ;
        RECT  18.330 3.055 18.525 3.725 ;
        RECT  17.990 3.055 18.330 3.865 ;
        RECT  17.800 1.280 18.140 1.850 ;
        RECT  16.890 2.080 18.100 2.420 ;
        RECT  16.835 2.080 16.890 3.340 ;
        RECT  16.660 1.505 16.835 3.340 ;
        RECT  16.605 1.505 16.660 2.310 ;
        RECT  16.550 2.975 16.660 3.340 ;
        RECT  16.165 1.505 16.605 1.735 ;
        RECT  15.450 2.975 16.550 3.205 ;
        RECT  15.920 2.130 16.260 2.470 ;
        RECT  15.930 1.055 16.165 1.735 ;
        RECT  15.800 1.055 15.930 1.580 ;
        RECT  13.495 2.185 15.920 2.415 ;
        RECT  14.415 1.055 15.800 1.285 ;
        RECT  15.340 2.975 15.450 3.340 ;
        RECT  15.110 2.975 15.340 3.725 ;
        RECT  14.120 3.495 15.110 3.725 ;
        RECT  14.075 1.000 14.415 1.340 ;
        RECT  13.835 3.495 14.120 4.040 ;
        RECT  13.780 3.700 13.835 4.040 ;
        RECT  13.275 0.810 13.615 1.150 ;
        RECT  13.325 1.385 13.495 3.165 ;
        RECT  13.265 1.385 13.325 3.260 ;
        RECT  12.045 0.865 13.275 1.095 ;
        RECT  12.995 1.385 13.265 1.770 ;
        RECT  12.985 2.915 13.265 3.260 ;
        RECT  12.690 2.220 13.030 2.560 ;
        RECT  11.380 1.385 12.995 1.615 ;
        RECT  11.300 2.915 12.985 3.145 ;
        RECT  12.145 2.220 12.690 2.450 ;
        RECT  11.915 1.980 12.145 2.450 ;
        RECT  11.815 0.675 12.045 1.095 ;
        RECT  11.720 1.980 11.915 2.210 ;
        RECT  10.740 0.675 11.815 0.905 ;
        RECT  11.380 1.870 11.720 2.210 ;
        RECT  11.040 1.160 11.380 1.615 ;
        RECT  10.960 2.915 11.300 3.440 ;
        RECT  10.655 2.310 11.050 2.650 ;
        RECT  10.655 0.675 10.740 1.600 ;
        RECT  10.510 0.675 10.655 3.100 ;
        RECT  10.425 1.370 10.510 3.100 ;
        RECT  9.260 1.370 10.425 1.600 ;
        RECT  9.345 2.870 10.425 3.100 ;
        RECT  8.855 2.270 10.190 2.610 ;
        RECT  9.115 2.870 9.345 3.265 ;
        RECT  8.920 0.700 9.260 1.600 ;
        RECT  8.745 3.035 9.115 3.265 ;
        RECT  8.700 3.520 9.040 4.010 ;
        RECT  8.765 0.700 8.920 1.040 ;
        RECT  8.455 2.230 8.855 2.610 ;
        RECT  6.155 3.520 8.700 3.750 ;
        RECT  8.295 1.715 8.455 3.265 ;
        RECT  8.225 0.960 8.295 3.265 ;
        RECT  8.065 0.960 8.225 1.945 ;
        RECT  6.785 3.035 8.225 3.265 ;
        RECT  7.955 0.960 8.065 1.300 ;
        RECT  7.645 2.400 7.930 2.740 ;
        RECT  7.415 1.450 7.645 2.740 ;
        RECT  5.655 1.450 7.415 1.680 ;
        RECT  6.555 2.010 6.785 3.265 ;
        RECT  6.445 2.010 6.555 2.350 ;
        RECT  5.925 2.020 6.155 4.235 ;
        RECT  5.705 2.020 5.925 2.360 ;
        RECT  5.275 4.005 5.925 4.235 ;
        RECT  5.475 3.000 5.690 3.720 ;
        RECT  5.475 1.000 5.655 1.680 ;
        RECT  5.460 1.000 5.475 3.720 ;
        RECT  5.315 1.000 5.460 3.230 ;
        RECT  5.245 1.450 5.315 3.230 ;
        RECT  4.935 3.950 5.275 4.290 ;
        RECT  4.645 3.135 4.985 3.570 ;
        RECT  4.350 4.005 4.935 4.235 ;
        RECT  4.510 0.730 4.850 1.070 ;
        RECT  2.205 3.135 4.645 3.365 ;
        RECT  2.215 0.840 4.510 1.070 ;
        RECT  4.120 3.675 4.350 4.235 ;
        RECT  2.560 3.675 4.120 3.905 ;
        RECT  3.430 1.330 3.770 1.670 ;
        RECT  2.300 1.405 3.430 1.635 ;
        RECT  2.330 3.675 2.560 4.105 ;
        RECT  2.300 2.490 2.505 2.905 ;
        RECT  0.520 3.875 2.330 4.105 ;
        RECT  2.070 1.405 2.300 2.905 ;
        RECT  1.985 0.630 2.215 1.070 ;
        RECT  1.840 2.675 2.070 2.905 ;
        RECT  1.790 0.630 1.985 0.860 ;
        RECT  1.610 2.675 1.840 3.620 ;
        RECT  1.500 3.280 1.610 3.620 ;
        RECT  0.410 1.270 0.520 1.610 ;
        RECT  0.410 2.960 0.520 4.105 ;
        RECT  0.290 1.270 0.410 4.105 ;
        RECT  0.180 1.270 0.290 3.300 ;
    END
END SDFFNSX4

MACRO SDFFNSX2
    CLASS CORE ;
    FOREIGN SDFFNSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.555 3.995 13.195 4.400 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 2.150 3.810 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.700 1.860 2.250 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.965 1.390 15.040 1.820 ;
        RECT  14.965 2.635 15.040 3.080 ;
        RECT  14.735 1.390 14.965 3.080 ;
        RECT  14.700 1.390 14.735 1.820 ;
        RECT  14.700 2.635 14.735 3.080 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.125 1.285 16.355 3.080 ;
        RECT  16.055 1.285 16.125 1.730 ;
        RECT  15.980 2.740 16.125 3.080 ;
        RECT  15.980 1.390 16.055 1.730 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.845 4.405 2.075 ;
        RECT  4.100 1.330 4.340 2.075 ;
        RECT  4.000 1.330 4.100 1.670 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.280 1.180 2.700 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.680 -0.400 16.500 0.400 ;
        RECT  15.340 -0.400 15.680 0.985 ;
        RECT  13.710 -0.400 15.340 0.400 ;
        RECT  13.370 -0.400 13.710 0.575 ;
        RECT  11.680 -0.400 13.370 0.400 ;
        RECT  11.340 -0.400 11.680 0.575 ;
        RECT  9.110 -0.400 11.340 0.400 ;
        RECT  8.880 -0.400 9.110 1.135 ;
        RECT  6.800 -0.400 8.880 0.400 ;
        RECT  6.460 -0.400 6.800 1.065 ;
        RECT  3.275 -0.400 6.460 0.400 ;
        RECT  2.935 -0.400 3.275 0.575 ;
        RECT  1.200 -0.400 2.935 0.400 ;
        RECT  0.860 -0.400 1.200 0.575 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.680 4.640 16.500 5.440 ;
        RECT  15.340 4.090 15.680 5.440 ;
        RECT  13.780 4.640 15.340 5.440 ;
        RECT  13.725 4.465 13.780 5.440 ;
        RECT  13.495 4.355 13.725 5.440 ;
        RECT  13.440 4.465 13.495 5.440 ;
        RECT  12.245 4.640 13.440 5.440 ;
        RECT  11.905 4.140 12.245 5.440 ;
        RECT  9.805 4.640 11.905 5.440 ;
        RECT  9.465 3.470 9.805 5.440 ;
        RECT  8.335 4.640 9.465 5.440 ;
        RECT  7.995 4.095 8.335 5.440 ;
        RECT  7.045 4.640 7.995 5.440 ;
        RECT  6.705 4.465 7.045 5.440 ;
        RECT  3.660 4.640 6.705 5.440 ;
        RECT  3.320 4.155 3.660 5.440 ;
        RECT  1.080 4.640 3.320 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.750 2.110 15.895 2.450 ;
        RECT  15.520 2.110 15.750 3.860 ;
        RECT  14.375 3.630 15.520 3.860 ;
        RECT  14.145 1.300 14.375 3.860 ;
        RECT  13.990 1.300 14.145 1.640 ;
        RECT  14.000 2.920 14.145 3.260 ;
        RECT  13.575 2.140 13.915 2.480 ;
        RECT  13.155 2.195 13.575 2.425 ;
        RECT  13.005 1.620 13.155 3.345 ;
        RECT  12.925 1.620 13.005 3.635 ;
        RECT  12.380 1.620 12.925 1.850 ;
        RECT  12.665 2.825 12.925 3.635 ;
        RECT  12.330 2.140 12.670 2.480 ;
        RECT  12.040 1.330 12.380 1.850 ;
        RECT  11.140 2.195 12.330 2.425 ;
        RECT  11.850 1.620 12.040 1.850 ;
        RECT  11.510 1.620 11.850 1.960 ;
        RECT  10.910 1.300 11.140 3.890 ;
        RECT  9.855 0.675 10.930 0.905 ;
        RECT  10.520 1.300 10.910 1.530 ;
        RECT  10.745 3.550 10.910 3.890 ;
        RECT  9.855 2.515 10.680 2.915 ;
        RECT  10.180 1.190 10.520 1.530 ;
        RECT  9.625 0.675 9.855 2.915 ;
        RECT  8.650 1.370 9.625 1.600 ;
        RECT  9.100 2.685 9.625 2.915 ;
        RECT  9.055 1.885 9.395 2.225 ;
        RECT  8.870 2.685 9.100 3.405 ;
        RECT  8.435 1.885 9.055 2.115 ;
        RECT  8.760 3.065 8.870 3.405 ;
        RECT  8.585 3.635 8.815 4.040 ;
        RECT  8.420 0.750 8.650 1.600 ;
        RECT  6.280 3.635 8.585 3.865 ;
        RECT  8.205 1.885 8.435 3.370 ;
        RECT  8.250 0.750 8.420 0.980 ;
        RECT  7.910 0.630 8.250 0.980 ;
        RECT  8.190 1.885 8.205 2.115 ;
        RECT  7.105 3.140 8.205 3.370 ;
        RECT  7.960 1.450 8.190 2.115 ;
        RECT  7.625 2.450 7.965 2.790 ;
        RECT  7.295 0.630 7.910 0.860 ;
        RECT  7.395 1.295 7.625 2.680 ;
        RECT  5.435 1.295 7.395 1.525 ;
        RECT  6.875 2.090 7.105 3.370 ;
        RECT  6.735 2.090 6.875 2.320 ;
        RECT  6.395 1.980 6.735 2.320 ;
        RECT  6.050 2.570 6.280 4.030 ;
        RECT  5.945 2.570 6.050 2.800 ;
        RECT  5.300 3.800 6.050 4.030 ;
        RECT  5.715 1.755 5.945 2.800 ;
        RECT  5.480 3.180 5.820 3.520 ;
        RECT  5.460 1.755 5.715 2.095 ;
        RECT  5.250 2.595 5.480 3.520 ;
        RECT  5.145 0.860 5.435 1.525 ;
        RECT  4.960 3.800 5.300 4.140 ;
        RECT  5.145 2.595 5.250 2.825 ;
        RECT  5.095 0.860 5.145 2.825 ;
        RECT  4.915 1.295 5.095 2.825 ;
        RECT  4.680 3.110 5.020 3.450 ;
        RECT  4.225 3.800 4.960 4.030 ;
        RECT  2.540 3.170 4.680 3.400 ;
        RECT  4.295 0.740 4.635 1.095 ;
        RECT  1.925 0.865 4.295 1.095 ;
        RECT  3.995 3.690 4.225 4.030 ;
        RECT  2.970 3.690 3.995 3.920 ;
        RECT  3.260 1.330 3.600 1.670 ;
        RECT  2.430 1.440 3.260 1.670 ;
        RECT  2.740 3.690 2.970 4.175 ;
        RECT  2.430 2.545 2.780 2.775 ;
        RECT  0.520 3.945 2.740 4.175 ;
        RECT  2.200 3.060 2.540 3.400 ;
        RECT  2.090 1.440 2.430 2.775 ;
        RECT  1.840 2.545 2.090 2.775 ;
        RECT  1.560 0.695 1.925 1.095 ;
        RECT  1.610 2.545 1.840 3.610 ;
        RECT  1.500 3.270 1.610 3.610 ;
        RECT  0.395 1.195 0.540 1.535 ;
        RECT  0.395 3.360 0.520 4.175 ;
        RECT  0.290 1.195 0.395 4.175 ;
        RECT  0.165 1.195 0.290 3.725 ;
    END
END SDFFNSX2

MACRO SDFFNSX1
    CLASS CORE ;
    FOREIGN SDFFNSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.985 3.770 13.270 4.110 ;
        RECT  12.755 3.770 12.985 4.315 ;
        RECT  12.680 3.770 12.755 4.060 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 2.150 3.810 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.470 1.700 1.870 2.250 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.965 0.860 15.015 3.755 ;
        RECT  14.890 0.860 14.965 3.850 ;
        RECT  14.785 0.860 14.890 4.085 ;
        RECT  14.300 0.860 14.785 1.090 ;
        RECT  14.735 3.525 14.785 4.085 ;
        RECT  14.660 3.620 14.735 4.085 ;
        RECT  14.360 3.855 14.660 4.085 ;
        RECT  14.020 3.855 14.360 4.195 ;
        RECT  13.960 0.750 14.300 1.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.640 3.095 15.660 3.435 ;
        RECT  15.320 1.210 15.640 3.435 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.330 4.405 2.075 ;
        RECT  4.100 1.330 4.175 1.820 ;
        RECT  3.960 1.330 4.100 1.670 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.685 2.280 1.180 2.700 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.020 -0.400 15.840 0.400 ;
        RECT  14.680 -0.400 15.020 0.575 ;
        RECT  13.500 -0.400 14.680 0.400 ;
        RECT  13.160 -0.400 13.500 0.575 ;
        RECT  11.680 -0.400 13.160 0.400 ;
        RECT  11.340 -0.400 11.680 0.575 ;
        RECT  9.110 -0.400 11.340 0.400 ;
        RECT  8.880 -0.400 9.110 1.100 ;
        RECT  6.800 -0.400 8.880 0.400 ;
        RECT  6.460 -0.400 6.800 1.065 ;
        RECT  3.275 -0.400 6.460 0.400 ;
        RECT  2.935 -0.400 3.275 0.575 ;
        RECT  1.200 -0.400 2.935 0.400 ;
        RECT  0.860 -0.400 1.200 0.575 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.150 4.640 15.840 5.440 ;
        RECT  14.715 4.465 15.150 5.440 ;
        RECT  13.600 4.640 14.715 5.440 ;
        RECT  13.260 4.465 13.600 5.440 ;
        RECT  12.320 4.640 13.260 5.440 ;
        RECT  11.980 4.140 12.320 5.440 ;
        RECT  9.825 4.640 11.980 5.440 ;
        RECT  9.485 3.635 9.825 5.440 ;
        RECT  8.335 4.640 9.485 5.440 ;
        RECT  7.995 4.095 8.335 5.440 ;
        RECT  7.045 4.640 7.995 5.440 ;
        RECT  6.705 4.465 7.045 5.440 ;
        RECT  3.660 4.640 6.705 5.440 ;
        RECT  3.320 4.155 3.660 5.440 ;
        RECT  1.080 4.640 3.320 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.325 1.600 14.555 3.145 ;
        RECT  14.300 1.600 14.325 1.830 ;
        RECT  14.020 2.805 14.325 3.145 ;
        RECT  13.960 1.490 14.300 1.830 ;
        RECT  13.600 2.140 13.940 2.480 ;
        RECT  13.080 2.195 13.600 2.425 ;
        RECT  12.850 1.620 13.080 3.400 ;
        RECT  12.380 1.620 12.850 1.850 ;
        RECT  12.690 3.060 12.850 3.400 ;
        RECT  12.280 2.380 12.620 2.720 ;
        RECT  12.040 1.190 12.380 1.850 ;
        RECT  11.140 2.435 12.280 2.665 ;
        RECT  11.850 1.620 12.040 1.850 ;
        RECT  11.510 1.620 11.850 1.960 ;
        RECT  10.910 1.545 11.140 3.890 ;
        RECT  9.855 0.675 10.930 0.905 ;
        RECT  10.520 1.545 10.910 1.775 ;
        RECT  10.765 3.550 10.910 3.890 ;
        RECT  9.855 2.515 10.680 2.915 ;
        RECT  10.290 1.190 10.520 1.775 ;
        RECT  10.180 1.190 10.290 1.530 ;
        RECT  9.625 0.675 9.855 2.915 ;
        RECT  8.650 1.370 9.625 1.600 ;
        RECT  9.100 2.685 9.625 2.915 ;
        RECT  8.435 1.835 9.395 2.065 ;
        RECT  8.870 2.685 9.100 3.405 ;
        RECT  8.760 3.065 8.870 3.405 ;
        RECT  8.585 3.635 8.815 4.040 ;
        RECT  8.420 0.695 8.650 1.600 ;
        RECT  6.280 3.635 8.585 3.865 ;
        RECT  8.205 1.835 8.435 3.370 ;
        RECT  7.650 0.695 8.420 0.925 ;
        RECT  8.190 1.835 8.205 2.065 ;
        RECT  7.105 3.140 8.205 3.370 ;
        RECT  7.960 1.420 8.190 2.065 ;
        RECT  7.735 2.355 7.965 2.740 ;
        RECT  7.625 2.355 7.735 2.585 ;
        RECT  7.295 0.675 7.650 0.925 ;
        RECT  7.395 1.295 7.625 2.585 ;
        RECT  5.435 1.295 7.395 1.525 ;
        RECT  6.875 2.060 7.105 3.370 ;
        RECT  6.735 2.060 6.875 2.290 ;
        RECT  6.395 1.950 6.735 2.290 ;
        RECT  6.050 2.570 6.280 4.085 ;
        RECT  5.945 2.570 6.050 2.800 ;
        RECT  5.295 3.855 6.050 4.085 ;
        RECT  5.715 1.805 5.945 2.800 ;
        RECT  5.480 3.180 5.820 3.520 ;
        RECT  5.460 1.805 5.715 2.035 ;
        RECT  5.250 2.595 5.480 3.425 ;
        RECT  5.145 0.860 5.435 1.525 ;
        RECT  4.955 3.800 5.295 4.140 ;
        RECT  5.145 2.595 5.250 2.825 ;
        RECT  5.095 0.860 5.145 2.825 ;
        RECT  4.915 1.295 5.095 2.825 ;
        RECT  4.680 3.110 5.020 3.450 ;
        RECT  4.345 3.800 4.955 4.030 ;
        RECT  2.540 3.165 4.680 3.395 ;
        RECT  4.295 0.740 4.635 1.080 ;
        RECT  4.115 3.690 4.345 4.030 ;
        RECT  1.900 0.850 4.295 1.080 ;
        RECT  2.970 3.690 4.115 3.920 ;
        RECT  3.260 1.330 3.600 1.670 ;
        RECT  2.375 1.385 3.260 1.615 ;
        RECT  2.740 3.690 2.970 4.175 ;
        RECT  2.440 2.490 2.780 2.830 ;
        RECT  0.520 3.945 2.740 4.175 ;
        RECT  2.200 3.060 2.540 3.400 ;
        RECT  2.375 2.490 2.440 2.775 ;
        RECT  2.145 1.385 2.375 2.775 ;
        RECT  1.840 2.545 2.145 2.775 ;
        RECT  1.560 0.640 1.900 1.080 ;
        RECT  1.610 2.545 1.840 3.610 ;
        RECT  1.500 3.270 1.610 3.610 ;
        RECT  0.395 1.195 0.540 1.535 ;
        RECT  0.395 3.360 0.520 4.175 ;
        RECT  0.290 1.195 0.395 4.175 ;
        RECT  0.165 1.195 0.290 3.725 ;
    END
END SDFFNSX1

MACRO SDFFNRXL
    CLASS CORE ;
    FOREIGN SDFFNRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 2.320 3.790 2.675 ;
        RECT  3.335 2.320 3.675 2.925 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 1.800 1.810 2.290 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.230 2.900 7.570 3.240 ;
        RECT  7.120 2.900 7.230 3.185 ;
        RECT  6.890 2.360 7.120 3.185 ;
        RECT  6.760 2.360 6.890 2.680 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.765 0.865 16.995 4.035 ;
        RECT  16.410 0.865 16.765 1.095 ;
        RECT  16.615 3.500 16.765 4.035 ;
        RECT  16.490 3.805 16.615 4.035 ;
        RECT  16.150 3.805 16.490 4.230 ;
        RECT  16.070 0.635 16.410 1.095 ;
        RECT  16.110 3.805 16.150 4.175 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.135 3.620 18.220 3.960 ;
        RECT  17.905 1.890 18.135 3.960 ;
        RECT  17.820 1.890 17.905 2.120 ;
        RECT  17.880 3.620 17.905 3.960 ;
        RECT  17.300 1.190 17.820 2.120 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.105 1.575 4.495 2.105 ;
        RECT  4.035 1.715 4.105 2.080 ;
        RECT  3.980 1.740 4.035 2.080 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.715 1.180 3.220 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.140 -0.400 18.480 0.400 ;
        RECT  16.800 -0.400 17.140 0.575 ;
        RECT  15.530 -0.400 16.800 0.400 ;
        RECT  15.190 -0.400 15.530 0.950 ;
        RECT  13.770 -0.400 15.190 0.400 ;
        RECT  13.430 -0.400 13.770 1.110 ;
        RECT  9.005 -0.400 13.430 0.400 ;
        RECT  10.535 1.205 10.875 1.760 ;
        RECT  9.300 1.205 10.535 1.435 ;
        RECT  9.005 1.205 9.300 1.580 ;
        RECT  8.960 -0.400 9.005 1.580 ;
        RECT  8.775 -0.400 8.960 1.525 ;
        RECT  6.990 -0.400 8.775 0.400 ;
        RECT  6.650 -0.400 6.990 0.960 ;
        RECT  3.300 -0.400 6.650 0.400 ;
        RECT  2.960 -0.400 3.300 0.575 ;
        RECT  1.210 -0.400 2.960 0.400 ;
        RECT  0.870 -0.400 1.210 0.575 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.450 4.640 18.480 5.440 ;
        RECT  17.110 4.465 17.450 5.440 ;
        RECT  15.730 4.640 17.110 5.440 ;
        RECT  15.390 4.110 15.730 5.440 ;
        RECT  13.705 4.640 15.390 5.440 ;
        RECT  13.365 4.080 13.705 5.440 ;
        RECT  11.370 4.640 13.365 5.440 ;
        RECT  10.430 4.080 11.370 5.440 ;
        RECT  7.300 4.640 10.430 5.440 ;
        RECT  6.960 4.465 7.300 5.440 ;
        RECT  3.730 4.640 6.960 5.440 ;
        RECT  3.390 4.080 3.730 5.440 ;
        RECT  0.760 4.640 3.390 5.440 ;
        RECT  0.420 4.465 0.760 5.440 ;
        RECT  0.000 4.640 0.420 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.380 1.380 16.490 3.160 ;
        RECT  16.150 1.380 16.380 3.350 ;
        RECT  15.970 1.380 16.150 1.850 ;
        RECT  16.040 2.820 16.150 3.350 ;
        RECT  15.625 1.880 15.670 2.220 ;
        RECT  15.615 1.865 15.625 2.220 ;
        RECT  15.115 1.865 15.615 2.245 ;
        RECT  14.885 1.865 15.115 3.850 ;
        RECT  14.675 1.865 14.885 2.095 ;
        RECT  14.410 3.620 14.885 3.850 ;
        RECT  14.445 0.915 14.675 2.095 ;
        RECT  14.310 3.005 14.650 3.390 ;
        RECT  14.285 0.915 14.445 1.825 ;
        RECT  14.070 3.620 14.410 3.960 ;
        RECT  13.175 3.160 14.310 3.390 ;
        RECT  13.875 1.595 14.285 1.825 ;
        RECT  13.875 2.240 13.930 2.580 ;
        RECT  13.645 1.595 13.875 2.580 ;
        RECT  13.590 2.240 13.645 2.580 ;
        RECT  12.995 1.425 13.175 3.405 ;
        RECT  12.995 4.000 13.000 4.340 ;
        RECT  12.945 1.425 12.995 4.340 ;
        RECT  12.230 1.425 12.945 1.655 ;
        RECT  12.765 3.160 12.945 4.340 ;
        RECT  12.660 4.000 12.765 4.340 ;
        RECT  12.255 2.390 12.595 2.730 ;
        RECT  12.170 0.630 12.510 0.970 ;
        RECT  11.575 2.445 12.255 2.675 ;
        RECT  11.945 1.290 12.230 1.655 ;
        RECT  11.575 0.685 12.170 0.915 ;
        RECT  11.890 1.290 11.945 1.630 ;
        RECT  11.345 0.675 11.575 3.465 ;
        RECT  9.955 0.675 11.345 0.915 ;
        RECT  10.790 3.075 11.345 3.465 ;
        RECT  9.615 2.140 11.030 2.480 ;
        RECT  10.495 2.810 10.550 3.150 ;
        RECT  10.265 2.810 10.495 3.825 ;
        RECT  10.210 2.810 10.265 3.150 ;
        RECT  10.135 3.595 10.265 3.825 ;
        RECT  9.905 3.595 10.135 4.365 ;
        RECT  9.670 0.675 9.955 0.905 ;
        RECT  7.765 4.135 9.905 4.365 ;
        RECT  9.330 0.635 9.670 0.975 ;
        RECT  9.385 1.825 9.615 3.690 ;
        RECT  8.350 1.825 9.385 2.055 ;
        RECT  9.080 3.460 9.385 3.690 ;
        RECT  8.740 3.460 9.080 3.800 ;
        RECT  8.730 2.440 9.070 2.780 ;
        RECT  8.125 2.495 8.730 2.725 ;
        RECT  8.350 1.100 8.360 1.440 ;
        RECT  8.120 1.100 8.350 2.055 ;
        RECT  8.125 3.485 8.345 3.870 ;
        RECT  8.005 2.435 8.125 3.870 ;
        RECT  8.020 1.100 8.120 1.885 ;
        RECT  6.540 1.655 8.020 1.885 ;
        RECT  7.895 2.435 8.005 3.715 ;
        RECT  7.890 2.435 7.895 2.665 ;
        RECT  7.555 2.115 7.890 2.665 ;
        RECT  7.535 3.945 7.765 4.365 ;
        RECT  7.535 0.770 7.760 1.110 ;
        RECT  7.550 2.115 7.555 2.455 ;
        RECT  7.420 0.770 7.535 1.420 ;
        RECT  6.645 3.945 7.535 4.175 ;
        RECT  7.305 0.825 7.420 1.420 ;
        RECT  5.500 1.190 7.305 1.420 ;
        RECT  6.435 2.935 6.645 4.355 ;
        RECT  6.200 1.655 6.540 2.080 ;
        RECT  6.415 2.395 6.435 4.355 ;
        RECT  6.205 2.395 6.415 3.165 ;
        RECT  5.570 4.125 6.415 4.355 ;
        RECT  5.875 2.395 6.205 2.625 ;
        RECT  6.175 1.655 6.200 2.025 ;
        RECT  5.915 3.460 6.100 3.800 ;
        RECT  5.760 2.935 5.915 3.800 ;
        RECT  5.810 1.915 5.875 2.625 ;
        RECT  5.645 1.890 5.810 2.625 ;
        RECT  5.685 2.935 5.760 3.745 ;
        RECT  5.335 2.935 5.685 3.165 ;
        RECT  5.470 1.890 5.645 2.230 ;
        RECT  5.230 4.070 5.570 4.410 ;
        RECT  5.165 0.980 5.500 1.420 ;
        RECT  5.165 2.545 5.335 3.165 ;
        RECT  4.275 4.125 5.230 4.355 ;
        RECT  4.880 3.460 5.220 3.800 ;
        RECT  5.160 0.980 5.165 3.165 ;
        RECT  5.105 1.190 5.160 3.165 ;
        RECT  4.935 1.190 5.105 2.775 ;
        RECT  4.740 3.460 4.880 3.690 ;
        RECT  4.510 3.160 4.740 3.690 ;
        RECT  4.570 0.960 4.660 1.300 ;
        RECT  4.320 0.865 4.570 1.300 ;
        RECT  2.710 3.160 4.510 3.390 ;
        RECT  2.155 0.865 4.320 1.095 ;
        RECT  4.045 3.620 4.275 4.355 ;
        RECT  3.155 3.620 4.045 3.850 ;
        RECT  3.170 1.615 3.510 1.955 ;
        RECT  2.430 1.670 3.170 1.900 ;
        RECT  2.925 3.620 3.155 4.225 ;
        RECT  1.395 3.995 2.925 4.225 ;
        RECT  2.370 3.050 2.710 3.390 ;
        RECT  2.375 1.450 2.430 1.900 ;
        RECT  2.375 2.480 2.380 2.820 ;
        RECT  2.145 1.450 2.375 2.820 ;
        RECT  1.940 0.685 2.155 1.095 ;
        RECT  2.090 1.450 2.145 1.790 ;
        RECT  2.040 2.480 2.145 2.820 ;
        RECT  1.955 2.590 2.040 2.820 ;
        RECT  1.955 3.340 2.010 3.680 ;
        RECT  1.725 2.590 1.955 3.680 ;
        RECT  1.925 0.630 1.940 1.095 ;
        RECT  1.600 0.630 1.925 0.970 ;
        RECT  1.670 3.340 1.725 3.680 ;
        RECT  1.165 3.745 1.395 4.225 ;
        RECT  0.540 3.745 1.165 3.975 ;
        RECT  0.485 1.220 0.540 1.560 ;
        RECT  0.395 3.530 0.540 3.975 ;
        RECT  0.395 1.195 0.485 1.560 ;
        RECT  0.165 1.195 0.395 3.975 ;
    END
END SDFFNRXL

MACRO SDFFNRX4
    CLASS CORE ;
    FOREIGN SDFFNRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.225 2.050 3.565 2.635 ;
        RECT  2.855 2.060 3.225 2.635 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.290 1.780 2.340 ;
        RECT  1.470 1.285 1.765 2.340 ;
        RECT  1.430 1.285 1.470 2.300 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.320 2.745 7.780 3.495 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.600 1.195 20.980 3.220 ;
        RECT  20.580 1.195 20.600 1.535 ;
        RECT  20.580 2.780 20.600 3.120 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.200 1.260 22.300 3.120 ;
        RECT  21.920 1.195 22.200 3.120 ;
        RECT  21.915 1.195 21.920 2.075 ;
        RECT  21.860 2.780 21.920 3.120 ;
        RECT  21.860 1.195 21.915 1.535 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 1.850 4.440 2.740 ;
        RECT  4.035 1.845 4.405 2.740 ;
        RECT  4.020 1.850 4.035 2.740 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.660 2.350 1.120 2.835 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.840 -0.400 23.100 0.400 ;
        RECT  22.500 -0.400 22.840 0.950 ;
        RECT  21.560 -0.400 22.500 0.400 ;
        RECT  21.220 -0.400 21.560 0.950 ;
        RECT  20.235 -0.400 21.220 0.400 ;
        RECT  19.895 -0.400 20.235 0.575 ;
        RECT  18.910 -0.400 19.895 0.400 ;
        RECT  18.570 -0.400 18.910 0.950 ;
        RECT  17.470 -0.400 18.570 0.400 ;
        RECT  17.130 -0.400 17.470 0.950 ;
        RECT  16.010 -0.400 17.130 0.400 ;
        RECT  15.670 -0.400 16.010 0.950 ;
        RECT  14.240 -0.400 15.670 0.400 ;
        RECT  13.900 -0.400 14.240 0.575 ;
        RECT  11.645 -0.400 13.900 0.400 ;
        RECT  11.415 -0.400 11.645 1.475 ;
        RECT  9.790 -0.400 11.415 0.400 ;
        RECT  11.230 1.245 11.415 1.475 ;
        RECT  9.450 -0.400 9.790 0.960 ;
        RECT  7.780 -0.400 9.450 0.400 ;
        RECT  7.440 -0.400 7.780 1.335 ;
        RECT  3.240 -0.400 7.440 0.400 ;
        RECT  2.900 -0.400 3.240 0.575 ;
        RECT  1.080 -0.400 2.900 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.840 4.640 23.100 5.440 ;
        RECT  22.500 4.040 22.840 5.440 ;
        RECT  21.560 4.640 22.500 5.440 ;
        RECT  21.220 4.040 21.560 5.440 ;
        RECT  20.235 4.640 21.220 5.440 ;
        RECT  19.895 4.465 20.235 5.440 ;
        RECT  18.710 4.640 19.895 5.440 ;
        RECT  18.370 3.055 18.710 5.440 ;
        RECT  16.110 4.640 18.370 5.440 ;
        RECT  15.770 4.080 16.110 5.440 ;
        RECT  13.630 4.640 15.770 5.440 ;
        RECT  13.290 3.675 13.630 5.440 ;
        RECT  10.780 4.640 13.290 5.440 ;
        RECT  10.440 3.920 10.780 5.440 ;
        RECT  7.120 4.640 10.440 5.440 ;
        RECT  6.780 4.465 7.120 5.440 ;
        RECT  3.880 4.640 6.780 5.440 ;
        RECT  3.540 4.080 3.880 5.440 ;
        RECT  0.850 4.640 3.540 5.440 ;
        RECT  0.510 4.465 0.850 5.440 ;
        RECT  0.000 4.640 0.510 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.605 2.030 22.835 3.750 ;
        RECT  20.275 3.520 22.605 3.750 ;
        RECT  20.045 1.395 20.275 3.750 ;
        RECT  19.590 1.395 20.045 1.730 ;
        RECT  19.430 3.265 20.045 3.495 ;
        RECT  18.810 2.100 19.750 2.440 ;
        RECT  19.250 1.390 19.590 1.730 ;
        RECT  19.090 2.975 19.430 3.785 ;
        RECT  19.240 1.395 19.250 1.675 ;
        RECT  18.190 2.155 18.810 2.385 ;
        RECT  17.960 0.720 18.190 2.690 ;
        RECT  17.850 0.720 17.960 1.475 ;
        RECT  17.430 2.460 17.960 2.690 ;
        RECT  16.750 1.245 17.850 1.475 ;
        RECT  17.355 1.725 17.710 2.065 ;
        RECT  17.200 2.460 17.430 3.835 ;
        RECT  16.770 1.725 17.355 2.105 ;
        RECT  17.090 2.985 17.200 3.835 ;
        RECT  15.500 3.605 17.090 3.835 ;
        RECT  15.765 1.875 16.770 2.105 ;
        RECT  16.520 0.700 16.750 1.475 ;
        RECT  16.410 0.700 16.520 1.040 ;
        RECT  15.535 1.495 15.765 3.365 ;
        RECT  13.195 1.495 15.535 1.735 ;
        RECT  14.905 3.135 15.535 3.365 ;
        RECT  15.270 3.605 15.500 4.250 ;
        RECT  14.765 2.425 15.105 2.820 ;
        RECT  13.660 0.955 15.020 1.185 ;
        RECT  14.905 3.750 14.960 4.090 ;
        RECT  14.675 3.135 14.905 4.090 ;
        RECT  12.735 2.425 14.765 2.655 ;
        RECT  12.995 3.135 14.675 3.365 ;
        RECT  14.620 3.750 14.675 4.090 ;
        RECT  13.430 0.635 13.660 1.185 ;
        RECT  12.220 0.635 13.430 0.865 ;
        RECT  12.965 1.095 13.195 1.735 ;
        RECT  12.765 3.135 12.995 3.855 ;
        RECT  12.550 1.095 12.965 1.325 ;
        RECT  12.350 3.625 12.765 3.855 ;
        RECT  12.505 1.720 12.735 2.655 ;
        RECT  12.010 3.625 12.350 3.990 ;
        RECT  11.990 0.635 12.220 3.145 ;
        RECT  10.765 1.715 11.990 1.975 ;
        RECT  11.705 2.915 11.990 3.145 ;
        RECT  10.175 2.205 11.760 2.435 ;
        RECT  11.540 2.915 11.705 3.945 ;
        RECT  11.315 2.915 11.540 4.000 ;
        RECT  11.200 3.660 11.315 4.000 ;
        RECT  10.805 2.840 10.970 3.180 ;
        RECT  10.575 2.840 10.805 3.660 ;
        RECT  10.535 0.675 10.765 1.975 ;
        RECT  10.045 3.430 10.575 3.660 ;
        RECT  10.040 0.675 10.535 0.905 ;
        RECT  9.945 1.565 10.175 3.145 ;
        RECT  9.815 3.430 10.045 4.365 ;
        RECT  9.230 1.565 9.945 1.795 ;
        RECT  9.500 2.915 9.945 3.145 ;
        RECT  7.665 4.135 9.815 4.365 ;
        RECT  9.160 2.915 9.500 3.870 ;
        RECT  9.130 2.100 9.470 2.440 ;
        RECT  8.890 1.430 9.230 1.795 ;
        RECT  8.315 2.155 9.130 2.385 ;
        RECT  6.760 1.565 8.890 1.795 ;
        RECT  8.315 3.560 8.370 3.900 ;
        RECT  8.085 2.025 8.315 3.900 ;
        RECT  7.570 2.025 8.085 2.255 ;
        RECT  8.030 3.560 8.085 3.900 ;
        RECT  7.435 3.945 7.665 4.365 ;
        RECT  6.465 3.945 7.435 4.175 ;
        RECT  6.905 2.320 6.960 2.660 ;
        RECT  5.625 0.825 6.950 1.055 ;
        RECT  6.760 2.245 6.905 2.660 ;
        RECT  6.620 1.565 6.760 2.660 ;
        RECT  6.530 1.565 6.620 2.475 ;
        RECT  6.235 3.035 6.465 4.345 ;
        RECT  6.120 3.035 6.235 3.265 ;
        RECT  4.365 4.115 6.235 4.345 ;
        RECT  5.890 1.980 6.120 3.265 ;
        RECT  5.660 3.500 5.920 3.840 ;
        RECT  5.840 1.980 5.890 2.210 ;
        RECT  5.500 1.870 5.840 2.210 ;
        RECT  5.430 2.465 5.660 3.840 ;
        RECT  5.400 0.825 5.625 1.415 ;
        RECT  5.065 2.465 5.430 2.695 ;
        RECT  5.395 0.825 5.400 1.470 ;
        RECT  5.065 1.130 5.395 1.470 ;
        RECT  5.025 3.430 5.200 3.770 ;
        RECT  5.060 1.130 5.065 2.695 ;
        RECT  4.835 1.185 5.060 2.695 ;
        RECT  4.795 3.135 5.025 3.770 ;
        RECT  2.760 3.135 4.795 3.365 ;
        RECT  4.260 0.865 4.600 1.250 ;
        RECT  4.135 3.615 4.365 4.345 ;
        RECT  2.615 0.865 4.260 1.095 ;
        RECT  3.240 3.615 4.135 3.845 ;
        RECT  3.185 1.330 3.525 1.670 ;
        RECT  3.010 3.615 3.240 4.235 ;
        RECT  2.475 1.440 3.185 1.670 ;
        RECT  0.520 4.005 3.010 4.235 ;
        RECT  2.475 3.135 2.760 3.600 ;
        RECT  2.385 0.680 2.615 1.095 ;
        RECT  2.410 1.440 2.475 2.845 ;
        RECT  2.420 3.260 2.475 3.600 ;
        RECT  2.145 1.360 2.410 2.845 ;
        RECT  1.540 0.680 2.385 0.910 ;
        RECT  2.070 1.360 2.145 1.700 ;
        RECT  2.105 2.615 2.145 2.845 ;
        RECT  1.875 2.615 2.105 3.650 ;
        RECT  1.840 3.420 1.875 3.650 ;
        RECT  1.500 3.420 1.840 3.760 ;
        RECT  0.465 1.220 0.520 1.560 ;
        RECT  0.405 3.180 0.520 4.235 ;
        RECT  0.405 1.215 0.465 1.560 ;
        RECT  0.290 1.215 0.405 4.235 ;
        RECT  0.175 1.215 0.290 3.520 ;
    END
END SDFFNRX4

MACRO SDFFNRX2
    CLASS CORE ;
    FOREIGN SDFFNRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.830 2.260 3.435 2.680 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.240 1.795 1.560 ;
        RECT  1.715 1.930 1.770 2.270 ;
        RECT  1.485 1.240 1.715 2.270 ;
        RECT  1.430 1.930 1.485 2.270 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.245 2.875 7.300 3.390 ;
        RECT  6.960 2.755 7.245 3.390 ;
        RECT  6.815 2.755 6.960 3.335 ;
        RECT  6.770 2.875 6.815 3.240 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.265 1.650 18.350 2.130 ;
        RECT  18.205 1.645 18.265 2.130 ;
        RECT  18.205 2.930 18.260 3.270 ;
        RECT  18.020 1.645 18.205 3.270 ;
        RECT  17.975 1.370 18.020 3.270 ;
        RECT  17.790 1.370 17.975 2.130 ;
        RECT  17.920 2.930 17.975 3.270 ;
        RECT  17.680 1.370 17.790 1.710 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.580 0.955 19.645 3.230 ;
        RECT  19.570 0.955 19.580 3.270 ;
        RECT  19.345 0.685 19.570 3.270 ;
        RECT  19.230 0.685 19.345 1.625 ;
        RECT  19.240 2.910 19.345 3.270 ;
        RECT  19.210 2.930 19.240 3.270 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.840 1.550 4.480 2.120 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.965 1.800 1.150 2.120 ;
        RECT  0.625 1.715 0.965 2.820 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.790 -0.400 19.800 0.400 ;
        RECT  18.450 -0.400 18.790 1.045 ;
        RECT  16.760 -0.400 18.450 0.400 ;
        RECT  16.420 -0.400 16.760 1.190 ;
        RECT  15.270 -0.400 16.420 0.400 ;
        RECT  14.930 -0.400 15.270 0.575 ;
        RECT  13.180 -0.400 14.930 0.400 ;
        RECT  12.840 -0.400 13.180 0.575 ;
        RECT  10.680 -0.400 12.840 0.400 ;
        RECT  10.340 -0.400 10.680 1.370 ;
        RECT  8.980 -0.400 10.340 0.400 ;
        RECT  8.640 -0.400 8.980 0.960 ;
        RECT  7.760 -0.400 8.640 0.440 ;
        RECT  7.335 -0.400 7.760 1.335 ;
        RECT  3.140 -0.400 7.335 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.080 -0.400 2.800 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.900 4.640 19.800 5.440 ;
        RECT  18.560 4.080 18.900 5.440 ;
        RECT  16.840 4.640 18.560 5.440 ;
        RECT  16.500 3.680 16.840 5.440 ;
        RECT  14.060 4.640 16.500 5.440 ;
        RECT  13.720 4.080 14.060 5.440 ;
        RECT  11.400 4.640 13.720 5.440 ;
        RECT  9.900 4.080 11.400 5.440 ;
        RECT  7.000 4.640 9.900 5.440 ;
        RECT  6.660 4.465 7.000 5.440 ;
        RECT  3.840 4.640 6.660 5.440 ;
        RECT  3.500 3.980 3.840 5.440 ;
        RECT  1.080 4.640 3.500 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.885 1.910 19.115 2.655 ;
        RECT  18.840 2.425 18.885 2.655 ;
        RECT  18.610 2.425 18.840 3.805 ;
        RECT  17.560 3.575 18.610 3.805 ;
        RECT  17.450 3.575 17.560 4.020 ;
        RECT  17.450 0.665 17.520 1.005 ;
        RECT  17.220 0.665 17.450 4.020 ;
        RECT  17.180 0.665 17.220 1.005 ;
        RECT  16.935 1.590 16.990 2.045 ;
        RECT  16.705 1.590 16.935 3.165 ;
        RECT  16.650 1.590 16.705 2.045 ;
        RECT  16.160 2.935 16.705 3.165 ;
        RECT  16.040 1.815 16.650 2.045 ;
        RECT  15.930 2.935 16.160 3.510 ;
        RECT  15.810 0.910 16.040 2.045 ;
        RECT  15.380 3.280 15.930 3.510 ;
        RECT  15.700 0.910 15.810 1.250 ;
        RECT  15.130 1.815 15.810 2.045 ;
        RECT  15.270 3.280 15.380 3.620 ;
        RECT  15.040 3.280 15.270 4.270 ;
        RECT  14.690 2.460 15.190 2.800 ;
        RECT  14.845 1.630 15.130 2.045 ;
        RECT  14.760 3.930 15.040 4.270 ;
        RECT  14.790 1.630 14.845 1.970 ;
        RECT  14.560 2.460 14.690 3.335 ;
        RECT  14.355 1.685 14.560 3.335 ;
        RECT  14.180 0.635 14.460 0.975 ;
        RECT  14.330 1.270 14.355 3.335 ;
        RECT  14.125 1.270 14.330 1.915 ;
        RECT  14.320 2.680 14.330 3.335 ;
        RECT  13.305 3.105 14.320 3.335 ;
        RECT  14.120 0.635 14.180 1.040 ;
        RECT  12.100 1.270 14.125 1.500 ;
        RECT  13.950 0.690 14.120 1.040 ;
        RECT  14.045 2.205 14.100 2.435 ;
        RECT  13.815 2.205 14.045 2.440 ;
        RECT  12.580 0.810 13.950 1.040 ;
        RECT  13.425 2.210 13.815 2.440 ;
        RECT  13.195 2.040 13.425 2.440 ;
        RECT  13.075 3.105 13.305 3.480 ;
        RECT  12.320 2.040 13.195 2.270 ;
        RECT  12.740 3.250 13.075 3.480 ;
        RECT  12.400 3.250 12.740 3.590 ;
        RECT  12.350 0.630 12.580 1.040 ;
        RECT  12.160 2.600 12.500 2.940 ;
        RECT  11.395 0.630 12.350 0.860 ;
        RECT  12.035 1.735 12.320 2.270 ;
        RECT  11.640 2.655 12.160 2.885 ;
        RECT  11.870 1.090 12.100 1.500 ;
        RECT  11.980 1.735 12.035 2.075 ;
        RECT  11.700 1.090 11.870 1.430 ;
        RECT  11.410 1.705 11.640 3.570 ;
        RECT  11.395 1.705 11.410 1.935 ;
        RECT  10.470 3.205 11.410 3.570 ;
        RECT  11.165 0.630 11.395 1.935 ;
        RECT  10.840 2.170 11.180 2.885 ;
        RECT  9.880 1.705 11.165 1.935 ;
        RECT  9.215 2.170 10.840 2.400 ;
        RECT  10.170 2.630 10.510 2.970 ;
        RECT  10.015 2.740 10.170 2.970 ;
        RECT  9.785 2.740 10.015 3.725 ;
        RECT  9.875 1.205 9.880 1.935 ;
        RECT  9.765 1.150 9.875 1.935 ;
        RECT  9.575 3.495 9.785 3.725 ;
        RECT  9.535 0.665 9.765 1.935 ;
        RECT  9.345 3.495 9.575 4.355 ;
        RECT  9.270 0.665 9.535 0.895 ;
        RECT  7.465 4.125 9.345 4.355 ;
        RECT  8.985 1.575 9.215 3.185 ;
        RECT  8.480 1.575 8.985 1.805 ;
        RECT  8.795 2.955 8.985 3.185 ;
        RECT  8.795 3.470 8.850 3.810 ;
        RECT  8.565 2.955 8.795 3.810 ;
        RECT  8.415 2.140 8.755 2.480 ;
        RECT  8.510 3.470 8.565 3.810 ;
        RECT  8.250 1.455 8.480 1.805 ;
        RECT  7.985 2.195 8.415 2.425 ;
        RECT  8.140 1.455 8.250 1.795 ;
        RECT  6.320 1.565 8.140 1.795 ;
        RECT  7.985 3.550 8.040 3.890 ;
        RECT  7.755 2.195 7.985 3.890 ;
        RECT  7.750 2.195 7.755 2.425 ;
        RECT  7.700 3.550 7.755 3.890 ;
        RECT  7.200 2.030 7.750 2.425 ;
        RECT  7.235 3.945 7.465 4.355 ;
        RECT  6.345 3.945 7.235 4.175 ;
        RECT  6.720 0.675 7.060 1.110 ;
        RECT  5.300 0.675 6.720 0.905 ;
        RECT  6.115 2.395 6.345 4.255 ;
        RECT  5.990 1.565 6.320 2.085 ;
        RECT  5.585 2.395 6.115 2.625 ;
        RECT  5.200 4.025 6.115 4.255 ;
        RECT  5.980 1.745 5.990 2.085 ;
        RECT  5.685 3.300 5.740 3.640 ;
        RECT  5.400 3.280 5.685 3.640 ;
        RECT  5.580 1.655 5.585 2.625 ;
        RECT  5.355 1.600 5.580 2.625 ;
        RECT  5.005 3.280 5.400 3.510 ;
        RECT  5.240 1.600 5.355 1.940 ;
        RECT  5.070 0.675 5.300 1.270 ;
        RECT  4.860 3.970 5.200 4.310 ;
        RECT  4.965 0.905 5.070 1.270 ;
        RECT  4.965 2.375 5.005 3.510 ;
        RECT  4.775 0.905 4.965 3.510 ;
        RECT  4.385 3.970 4.860 4.200 ;
        RECT  4.735 0.905 4.775 2.605 ;
        RECT  4.205 2.850 4.545 3.190 ;
        RECT  4.160 0.865 4.500 1.285 ;
        RECT  4.155 3.450 4.385 4.200 ;
        RECT  2.475 2.935 4.205 3.165 ;
        RECT  2.565 0.865 4.160 1.095 ;
        RECT  2.515 3.450 4.155 3.680 ;
        RECT  3.020 1.635 3.360 1.975 ;
        RECT  2.410 1.690 3.020 1.920 ;
        RECT  2.335 0.665 2.565 1.095 ;
        RECT  2.285 3.450 2.515 4.235 ;
        RECT  2.230 1.460 2.410 2.070 ;
        RECT  1.785 0.665 2.335 0.895 ;
        RECT  0.520 4.005 2.285 4.235 ;
        RECT  2.070 1.460 2.230 2.740 ;
        RECT  2.065 1.840 2.070 2.740 ;
        RECT  2.000 1.840 2.065 3.180 ;
        RECT  1.880 2.505 2.000 3.180 ;
        RECT  1.835 2.505 1.880 3.770 ;
        RECT  1.650 2.840 1.835 3.770 ;
        RECT  1.440 0.665 1.785 0.960 ;
        RECT  1.540 3.430 1.650 3.770 ;
        RECT  0.395 1.100 0.520 1.440 ;
        RECT  0.395 3.630 0.520 4.235 ;
        RECT  0.165 1.100 0.395 4.235 ;
    END
END SDFFNRX2

MACRO SDFFNRX1
    CLASS CORE ;
    FOREIGN SDFFNRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNRXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 2.350 3.820 2.860 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.760 1.810 2.220 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.165 3.340 7.795 3.570 ;
        RECT  6.935 2.390 7.165 3.570 ;
        RECT  6.770 2.390 6.935 2.650 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.020 0.860 17.050 3.295 ;
        RECT  16.820 0.860 17.020 3.780 ;
        RECT  16.640 0.860 16.820 1.285 ;
        RECT  16.715 3.065 16.820 3.780 ;
        RECT  16.380 3.525 16.715 3.780 ;
        RECT  15.940 0.860 16.640 1.090 ;
        RECT  16.150 3.525 16.380 3.990 ;
        RECT  16.000 3.650 16.150 3.990 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.640 1.270 17.655 3.660 ;
        RECT  17.395 1.270 17.640 3.935 ;
        RECT  17.375 1.270 17.395 1.845 ;
        RECT  17.300 3.125 17.395 3.935 ;
        RECT  17.300 1.355 17.375 1.845 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 1.600 4.420 2.120 ;
        RECT  3.940 1.615 4.020 2.120 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.670 1.180 3.230 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.560 -0.400 17.820 0.400 ;
        RECT  17.220 -0.400 17.560 0.575 ;
        RECT  14.890 -0.400 17.220 0.400 ;
        RECT  14.550 -0.400 14.890 0.575 ;
        RECT  13.370 -0.400 14.550 0.400 ;
        RECT  13.030 -0.400 13.370 0.575 ;
        RECT  9.005 -0.400 13.030 0.400 ;
        RECT  10.780 1.440 10.890 1.780 ;
        RECT  10.550 1.205 10.780 1.780 ;
        RECT  9.300 1.205 10.550 1.435 ;
        RECT  9.005 1.205 9.300 1.525 ;
        RECT  8.775 -0.400 9.005 1.525 ;
        RECT  6.990 -0.400 8.775 0.400 ;
        RECT  6.650 -0.400 6.990 0.960 ;
        RECT  3.200 -0.400 6.650 0.400 ;
        RECT  2.860 -0.400 3.200 0.575 ;
        RECT  0.540 -0.400 2.860 0.400 ;
        RECT  0.200 -0.400 0.540 0.575 ;
        RECT  0.000 -0.400 0.200 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.550 4.640 17.820 5.440 ;
        RECT  17.110 4.465 17.550 5.440 ;
        RECT  15.620 4.640 17.110 5.440 ;
        RECT  15.280 3.620 15.620 5.440 ;
        RECT  13.640 4.640 15.280 5.440 ;
        RECT  13.300 4.070 13.640 5.440 ;
        RECT  11.370 4.640 13.300 5.440 ;
        RECT  10.430 4.070 11.370 5.440 ;
        RECT  7.300 4.640 10.430 5.440 ;
        RECT  6.960 4.465 7.300 5.440 ;
        RECT  3.730 4.640 6.960 5.440 ;
        RECT  3.390 4.080 3.730 5.440 ;
        RECT  1.130 4.640 3.390 5.440 ;
        RECT  0.790 4.465 1.130 5.440 ;
        RECT  0.000 4.640 0.790 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.365 2.150 16.420 2.490 ;
        RECT  16.230 2.145 16.365 2.490 ;
        RECT  15.935 2.145 16.230 3.110 ;
        RECT  15.890 1.320 15.935 3.110 ;
        RECT  15.705 1.320 15.890 2.375 ;
        RECT  15.440 1.320 15.705 1.550 ;
        RECT  15.245 1.825 15.475 3.295 ;
        RECT  15.100 1.210 15.440 1.550 ;
        RECT  14.810 1.825 15.245 2.055 ;
        RECT  14.340 3.065 15.245 3.295 ;
        RECT  14.580 1.595 14.810 2.055 ;
        RECT  14.130 1.595 14.580 1.825 ;
        RECT  14.010 2.140 14.350 2.480 ;
        RECT  14.110 3.065 14.340 3.815 ;
        RECT  13.790 0.680 14.130 1.825 ;
        RECT  14.000 3.475 14.110 3.815 ;
        RECT  12.830 2.245 14.010 2.475 ;
        RECT  13.450 1.595 13.790 1.825 ;
        RECT  13.110 1.595 13.450 2.015 ;
        RECT  12.830 4.000 12.940 4.340 ;
        RECT  12.600 2.020 12.830 4.340 ;
        RECT  12.155 2.020 12.600 2.250 ;
        RECT  12.190 0.665 12.530 1.005 ;
        RECT  12.120 2.500 12.230 2.840 ;
        RECT  12.155 1.310 12.210 1.650 ;
        RECT  11.575 0.675 12.190 0.905 ;
        RECT  11.925 1.310 12.155 2.250 ;
        RECT  11.890 2.500 12.120 3.330 ;
        RECT  11.870 1.310 11.925 1.650 ;
        RECT  11.575 3.100 11.890 3.330 ;
        RECT  11.345 0.675 11.575 3.330 ;
        RECT  9.575 0.675 11.345 0.905 ;
        RECT  10.955 3.100 11.345 3.330 ;
        RECT  10.690 2.020 11.030 2.410 ;
        RECT  10.725 3.100 10.955 3.575 ;
        RECT  9.615 2.180 10.690 2.410 ;
        RECT  10.265 2.705 10.495 3.825 ;
        RECT  10.135 3.595 10.265 3.825 ;
        RECT  9.905 3.595 10.135 4.365 ;
        RECT  7.760 4.135 9.905 4.365 ;
        RECT  9.385 1.825 9.615 3.385 ;
        RECT  9.235 0.635 9.575 0.975 ;
        RECT  8.485 1.825 9.385 2.055 ;
        RECT  9.080 3.155 9.385 3.385 ;
        RECT  8.850 3.155 9.080 3.820 ;
        RECT  8.730 2.440 9.070 2.780 ;
        RECT  8.740 3.480 8.850 3.820 ;
        RECT  8.325 2.495 8.730 2.725 ;
        RECT  8.255 1.115 8.485 2.055 ;
        RECT  8.325 3.480 8.380 3.820 ;
        RECT  8.095 2.435 8.325 3.820 ;
        RECT  8.075 1.115 8.255 1.885 ;
        RECT  7.890 2.435 8.095 2.665 ;
        RECT  8.040 3.480 8.095 3.820 ;
        RECT  6.540 1.655 8.075 1.885 ;
        RECT  7.525 2.120 7.890 2.665 ;
        RECT  7.535 0.770 7.830 1.110 ;
        RECT  7.530 3.945 7.760 4.365 ;
        RECT  7.305 0.770 7.535 1.420 ;
        RECT  6.645 3.945 7.530 4.175 ;
        RECT  5.500 1.190 7.305 1.420 ;
        RECT  6.435 2.935 6.645 4.320 ;
        RECT  6.200 1.655 6.540 2.080 ;
        RECT  6.415 2.395 6.435 4.320 ;
        RECT  6.205 2.395 6.415 3.165 ;
        RECT  4.275 4.090 6.415 4.320 ;
        RECT  5.875 2.395 6.205 2.625 ;
        RECT  5.745 3.480 6.080 3.840 ;
        RECT  5.645 1.940 5.875 2.625 ;
        RECT  5.515 2.855 5.745 3.840 ;
        RECT  5.480 1.940 5.645 2.280 ;
        RECT  5.340 2.855 5.515 3.085 ;
        RECT  5.165 1.160 5.500 1.500 ;
        RECT  5.165 2.590 5.340 3.085 ;
        RECT  4.910 3.435 5.250 3.800 ;
        RECT  5.110 1.160 5.165 3.085 ;
        RECT  4.935 1.160 5.110 2.820 ;
        RECT  4.795 3.435 4.910 3.665 ;
        RECT  4.565 3.100 4.795 3.665 ;
        RECT  2.730 3.100 4.565 3.330 ;
        RECT  4.220 0.865 4.560 1.250 ;
        RECT  4.045 3.620 4.275 4.320 ;
        RECT  2.155 0.865 4.220 1.095 ;
        RECT  3.120 3.620 4.045 3.850 ;
        RECT  3.170 1.330 3.510 1.670 ;
        RECT  2.430 1.385 3.170 1.615 ;
        RECT  2.890 3.620 3.120 3.975 ;
        RECT  0.550 3.745 2.890 3.975 ;
        RECT  2.390 3.045 2.730 3.385 ;
        RECT  2.375 2.460 2.580 2.800 ;
        RECT  2.375 1.385 2.430 1.750 ;
        RECT  2.240 1.385 2.375 2.800 ;
        RECT  2.145 1.385 2.240 2.745 ;
        RECT  1.925 0.665 2.155 1.095 ;
        RECT  2.090 1.385 2.145 1.750 ;
        RECT  1.990 2.515 2.145 2.745 ;
        RECT  1.760 2.515 1.990 3.240 ;
        RECT  1.500 0.665 1.925 0.895 ;
        RECT  1.650 2.900 1.760 3.240 ;
        RECT  0.395 3.520 0.550 3.975 ;
        RECT  0.395 1.350 0.540 1.690 ;
        RECT  0.165 1.350 0.395 3.975 ;
    END
END SDFFNRX1

MACRO SDFFNXL
    CLASS CORE ;
    FOREIGN SDFFNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 1.820 3.160 2.100 ;
        RECT  2.365 1.730 2.695 2.100 ;
        RECT  2.310 1.730 2.365 1.960 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.665 2.600 4.005 2.940 ;
        RECT  3.180 2.655 3.665 2.885 ;
        RECT  2.950 2.380 3.180 2.885 ;
        RECT  2.120 2.380 2.950 2.660 ;
        RECT  1.990 2.405 2.120 2.635 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.000 3.515 13.340 3.855 ;
        RECT  12.985 1.225 13.020 1.565 ;
        RECT  12.985 3.515 13.000 3.755 ;
        RECT  12.755 1.225 12.985 3.745 ;
        RECT  12.680 1.225 12.755 1.565 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.750 0.630 12.090 1.045 ;
        RECT  11.715 2.045 11.905 3.440 ;
        RECT  11.650 0.815 11.750 1.045 ;
        RECT  11.675 2.045 11.715 3.550 ;
        RECT  11.650 2.045 11.675 2.275 ;
        RECT  11.375 3.210 11.675 3.550 ;
        RECT  11.420 0.815 11.650 2.275 ;
        RECT  10.775 1.285 11.420 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 1.845 4.405 2.075 ;
        RECT  3.960 1.405 4.245 2.075 ;
        RECT  3.905 1.405 3.960 1.745 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.255 1.180 2.660 ;
        RECT  0.800 2.200 0.875 2.660 ;
        RECT  0.645 2.200 0.800 2.655 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.915 -0.400 13.860 0.400 ;
        RECT  12.575 -0.400 12.915 0.575 ;
        RECT  11.330 -0.400 12.575 0.400 ;
        RECT  10.990 -0.400 11.330 0.575 ;
        RECT  8.890 -0.400 10.990 0.400 ;
        RECT  8.550 -0.400 8.890 1.510 ;
        RECT  6.535 -0.400 8.550 0.400 ;
        RECT  6.305 -0.400 6.535 1.150 ;
        RECT  3.070 -0.400 6.305 0.400 ;
        RECT  2.730 -0.400 3.070 0.575 ;
        RECT  1.140 -0.400 2.730 0.400 ;
        RECT  1.140 1.290 1.320 1.630 ;
        RECT  0.980 -0.400 1.140 1.630 ;
        RECT  0.910 -0.400 0.980 1.575 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.515 4.640 13.860 5.440 ;
        RECT  12.175 4.410 12.515 5.440 ;
        RECT  10.915 4.640 12.175 5.440 ;
        RECT  10.575 4.465 10.915 5.440 ;
        RECT  8.215 4.640 10.575 5.440 ;
        RECT  6.935 4.465 8.215 5.440 ;
        RECT  4.005 4.640 6.935 5.440 ;
        RECT  3.665 4.410 4.005 5.440 ;
        RECT  0.940 4.640 3.665 5.440 ;
        RECT  0.530 4.465 0.940 5.440 ;
        RECT  0.000 4.640 0.530 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.220 1.415 12.450 4.180 ;
        RECT  11.880 1.360 12.220 1.700 ;
        RECT  11.735 3.950 12.220 4.180 ;
        RECT  11.505 3.950 11.735 4.350 ;
        RECT  11.285 4.005 11.505 4.350 ;
        RECT  11.180 2.615 11.435 2.955 ;
        RECT  10.545 4.005 11.285 4.235 ;
        RECT  11.095 2.260 11.180 2.955 ;
        RECT  10.950 2.260 11.095 2.845 ;
        RECT  10.170 2.260 10.950 2.490 ;
        RECT  9.415 0.795 10.570 1.025 ;
        RECT  10.315 2.745 10.545 4.235 ;
        RECT  10.205 2.745 10.315 3.085 ;
        RECT  9.880 1.310 10.170 2.490 ;
        RECT  9.830 1.310 9.880 4.150 ;
        RECT  9.755 2.260 9.830 4.150 ;
        RECT  9.650 2.260 9.755 4.260 ;
        RECT  9.415 3.920 9.650 4.260 ;
        RECT  9.305 0.795 9.415 3.260 ;
        RECT  9.185 0.795 9.305 3.615 ;
        RECT  8.090 1.740 9.185 1.970 ;
        RECT  9.075 2.920 9.185 3.615 ;
        RECT  8.910 3.385 9.075 3.615 ;
        RECT  8.615 2.200 8.955 2.540 ;
        RECT  8.680 3.385 8.910 4.235 ;
        RECT  6.325 4.005 8.680 4.235 ;
        RECT  8.440 2.310 8.615 2.540 ;
        RECT  8.210 2.310 8.440 3.775 ;
        RECT  7.300 3.545 8.210 3.775 ;
        RECT  7.875 1.170 8.090 1.970 ;
        RECT  7.750 1.170 7.875 3.120 ;
        RECT  7.745 1.225 7.750 3.120 ;
        RECT  7.645 1.740 7.745 3.120 ;
        RECT  7.535 2.780 7.645 3.120 ;
        RECT  7.300 0.810 7.390 1.150 ;
        RECT  7.070 0.810 7.300 3.775 ;
        RECT  7.050 0.810 7.070 1.150 ;
        RECT  6.760 2.275 7.070 2.505 ;
        RECT  6.500 1.550 6.840 1.890 ;
        RECT  6.420 2.220 6.760 2.560 ;
        RECT  6.015 1.605 6.500 1.835 ;
        RECT  6.270 3.780 6.325 4.235 ;
        RECT  6.040 3.715 6.270 4.235 ;
        RECT  5.985 3.715 6.040 4.120 ;
        RECT  5.890 0.795 6.015 1.835 ;
        RECT  5.430 3.715 5.985 3.945 ;
        RECT  5.660 0.795 5.890 3.480 ;
        RECT  4.890 0.795 5.660 1.025 ;
        RECT  4.900 4.180 5.460 4.410 ;
        RECT  5.200 1.760 5.430 3.945 ;
        RECT  4.955 1.760 5.200 1.990 ;
        RECT  4.630 3.320 4.970 3.660 ;
        RECT  4.725 1.390 4.955 1.990 ;
        RECT  4.670 3.920 4.900 4.410 ;
        RECT  3.435 3.920 4.670 4.150 ;
        RECT  2.975 3.430 4.630 3.660 ;
        RECT  4.090 0.750 4.430 1.090 ;
        RECT  2.485 0.810 4.090 1.040 ;
        RECT  3.195 1.345 3.460 1.575 ;
        RECT  3.205 3.920 3.435 4.410 ;
        RECT  1.895 4.180 3.205 4.410 ;
        RECT  2.965 1.270 3.195 1.575 ;
        RECT  2.745 3.430 2.975 3.930 ;
        RECT  2.065 1.270 2.965 1.500 ;
        RECT  2.150 3.700 2.745 3.930 ;
        RECT  2.255 0.645 2.485 1.040 ;
        RECT  2.145 3.040 2.485 3.380 ;
        RECT  1.370 0.645 2.255 0.875 ;
        RECT  1.860 3.040 2.145 3.270 ;
        RECT  1.835 1.270 2.065 2.150 ;
        RECT  1.665 3.605 1.895 4.410 ;
        RECT  1.750 2.905 1.860 3.270 ;
        RECT  1.750 1.920 1.835 2.150 ;
        RECT  1.520 1.920 1.750 3.270 ;
        RECT  0.540 3.605 1.665 3.835 ;
        RECT  0.380 2.995 0.540 3.835 ;
        RECT  0.380 1.430 0.520 1.770 ;
        RECT  0.310 1.430 0.380 3.835 ;
        RECT  0.200 1.430 0.310 3.335 ;
        RECT  0.180 1.430 0.200 3.225 ;
        RECT  0.150 1.485 0.180 3.225 ;
    END
END SDFFNXL

MACRO SDFFNX4
    CLASS CORE ;
    FOREIGN SDFFNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.790 1.820 3.320 2.240 ;
        RECT  2.780 1.820 2.790 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 2.545 3.870 2.775 ;
        RECT  2.245 2.380 2.500 2.775 ;
        RECT  2.010 2.380 2.245 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 1.820 17.680 3.220 ;
        RECT  17.300 1.460 17.605 3.220 ;
        RECT  17.265 1.460 17.300 1.845 ;
        RECT  17.295 2.635 17.300 3.110 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.325 1.820 16.360 3.220 ;
        RECT  15.985 1.460 16.325 3.220 ;
        RECT  15.980 1.820 15.985 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.405 4.405 2.635 ;
        RECT  4.380 1.550 4.385 2.635 ;
        RECT  4.150 1.495 4.380 2.635 ;
        RECT  4.040 1.495 4.150 1.835 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 2.200 1.105 2.635 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 -0.400 18.480 0.400 ;
        RECT  17.905 -0.400 18.245 1.090 ;
        RECT  16.965 -0.400 17.905 0.400 ;
        RECT  16.625 -0.400 16.965 1.090 ;
        RECT  15.645 -0.400 16.625 0.400 ;
        RECT  15.305 -0.400 15.645 0.575 ;
        RECT  14.225 -0.400 15.305 0.400 ;
        RECT  13.995 -0.400 14.225 1.310 ;
        RECT  11.585 -0.400 13.995 0.400 ;
        RECT  11.355 -0.400 11.585 1.335 ;
        RECT  9.025 -0.400 11.355 0.400 ;
        RECT  8.795 -0.400 9.025 1.370 ;
        RECT  6.740 -0.400 8.795 0.400 ;
        RECT  6.400 -0.400 6.740 1.270 ;
        RECT  3.220 -0.400 6.400 0.400 ;
        RECT  2.880 -0.400 3.220 0.575 ;
        RECT  1.290 -0.400 2.880 0.400 ;
        RECT  1.290 1.445 1.320 1.785 ;
        RECT  0.980 -0.400 1.290 1.785 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.275 4.640 18.480 5.440 ;
        RECT  17.935 4.090 18.275 5.440 ;
        RECT  16.970 4.640 17.935 5.440 ;
        RECT  16.630 4.090 16.970 5.440 ;
        RECT  15.690 4.640 16.630 5.440 ;
        RECT  15.350 4.090 15.690 5.440 ;
        RECT  14.250 4.640 15.350 5.440 ;
        RECT  13.860 4.465 14.250 5.440 ;
        RECT  11.775 4.640 13.860 5.440 ;
        RECT  11.435 4.005 11.775 5.440 ;
        RECT  9.150 4.640 11.435 5.440 ;
        RECT  8.810 4.465 9.150 5.440 ;
        RECT  6.980 4.640 8.810 5.440 ;
        RECT  6.640 4.465 6.980 5.440 ;
        RECT  1.380 4.640 6.640 5.440 ;
        RECT  1.040 4.465 1.380 5.440 ;
        RECT  0.000 4.640 1.040 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.910 2.055 18.140 3.860 ;
        RECT  14.925 3.630 17.910 3.860 ;
        RECT  15.520 1.285 15.750 3.020 ;
        RECT  15.000 1.285 15.520 1.570 ;
        RECT  14.925 2.700 15.520 3.020 ;
        RECT  14.475 2.040 15.285 2.380 ;
        RECT  14.660 1.230 15.000 1.570 ;
        RECT  14.585 2.700 14.925 3.865 ;
        RECT  14.015 2.700 14.585 2.930 ;
        RECT  13.755 2.095 14.475 2.325 ;
        RECT  13.675 2.645 14.015 2.985 ;
        RECT  13.525 0.970 13.755 2.325 ;
        RECT  12.920 0.970 13.525 1.250 ;
        RECT  13.170 2.095 13.525 2.325 ;
        RECT  12.690 1.550 13.290 1.780 ;
        RECT  13.060 2.095 13.170 3.780 ;
        RECT  12.940 2.095 13.060 4.070 ;
        RECT  12.720 3.260 12.940 4.070 ;
        RECT  12.580 0.965 12.920 1.305 ;
        RECT  10.490 3.450 12.720 3.680 ;
        RECT  12.635 1.550 12.690 2.935 ;
        RECT  12.460 1.550 12.635 2.970 ;
        RECT  12.230 1.075 12.580 1.305 ;
        RECT  12.350 2.595 12.460 2.970 ;
        RECT  12.185 2.740 12.350 2.970 ;
        RECT  12.000 1.075 12.230 1.805 ;
        RECT  11.955 2.740 12.185 3.040 ;
        RECT  10.960 1.575 12.000 1.805 ;
        RECT  10.730 2.810 11.955 3.040 ;
        RECT  11.660 2.235 11.715 2.575 ;
        RECT  11.375 2.035 11.660 2.575 ;
        RECT  9.450 2.035 11.375 2.265 ;
        RECT  10.730 1.250 10.960 1.805 ;
        RECT  10.360 1.250 10.730 1.480 ;
        RECT  10.445 2.595 10.730 3.040 ;
        RECT  10.150 3.450 10.490 4.260 ;
        RECT  10.390 2.595 10.445 3.000 ;
        RECT  8.640 2.650 10.390 3.000 ;
        RECT  10.020 1.140 10.360 1.480 ;
        RECT  9.395 2.035 9.450 2.400 ;
        RECT  9.165 1.600 9.395 2.400 ;
        RECT  8.565 1.600 9.165 1.830 ;
        RECT  9.110 2.060 9.165 2.400 ;
        RECT  8.410 2.650 8.640 4.235 ;
        RECT  8.335 0.630 8.565 1.830 ;
        RECT  8.255 2.650 8.410 3.655 ;
        RECT  5.540 4.005 8.410 4.235 ;
        RECT  7.460 0.630 8.335 0.860 ;
        RECT  8.105 2.650 8.255 2.880 ;
        RECT  8.200 3.315 8.255 3.655 ;
        RECT  7.875 1.175 8.105 2.880 ;
        RECT  7.445 3.320 7.785 3.660 ;
        RECT  7.435 0.630 7.460 1.485 ;
        RECT  7.440 3.320 7.445 3.605 ;
        RECT  7.435 2.575 7.440 3.605 ;
        RECT  7.230 0.630 7.435 3.605 ;
        RECT  7.210 1.145 7.230 3.605 ;
        RECT  7.205 1.145 7.210 3.550 ;
        RECT  7.120 1.145 7.205 1.485 ;
        RECT  6.815 2.575 7.205 2.805 ;
        RECT  5.810 1.905 6.975 2.135 ;
        RECT  6.475 2.520 6.815 2.860 ;
        RECT  5.580 0.685 5.810 3.490 ;
        RECT  5.040 0.685 5.580 0.915 ;
        RECT  5.350 3.720 5.540 4.235 ;
        RECT  5.310 2.820 5.350 4.235 ;
        RECT  5.120 2.820 5.310 3.950 ;
        RECT  4.995 2.820 5.120 3.050 ;
        RECT  1.840 4.180 5.080 4.410 ;
        RECT  4.765 1.390 4.995 3.050 ;
        RECT  3.860 3.315 4.890 3.545 ;
        RECT  4.525 0.670 4.580 1.010 ;
        RECT  4.240 0.670 4.525 1.035 ;
        RECT  2.650 0.805 4.240 1.035 ;
        RECT  3.630 3.315 3.860 3.930 ;
        RECT  2.155 1.335 3.630 1.565 ;
        RECT  2.070 3.700 3.630 3.930 ;
        RECT  2.420 0.645 2.650 1.035 ;
        RECT  1.940 3.095 2.650 3.325 ;
        RECT  1.520 0.645 2.420 0.875 ;
        RECT  1.925 1.335 2.155 2.150 ;
        RECT  1.780 2.905 1.940 3.325 ;
        RECT  1.780 1.920 1.925 2.150 ;
        RECT  1.610 4.005 1.840 4.410 ;
        RECT  1.550 1.920 1.780 3.325 ;
        RECT  0.620 4.005 1.610 4.235 ;
        RECT  0.350 2.880 0.620 4.235 ;
        RECT  0.350 0.985 0.600 1.795 ;
        RECT  0.280 0.985 0.350 4.235 ;
        RECT  0.260 0.985 0.280 3.255 ;
        RECT  0.120 1.275 0.260 3.255 ;
    END
END SDFFNX4

MACRO SDFFNX2
    CLASS CORE ;
    FOREIGN SDFFNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.980 1.820 3.160 2.100 ;
        RECT  2.470 1.730 2.980 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.055 2.695 4.165 3.035 ;
        RECT  3.825 2.405 4.055 3.035 ;
        RECT  3.745 2.405 3.825 2.660 ;
        RECT  2.500 2.405 3.745 2.635 ;
        RECT  2.050 2.380 2.500 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.395 1.355 15.625 3.170 ;
        RECT  15.320 1.355 15.395 1.845 ;
        RECT  15.340 2.940 15.395 3.195 ;
        RECT  15.000 2.940 15.340 3.750 ;
        RECT  15.220 1.355 15.320 1.695 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.860 0.700 14.200 1.080 ;
        RECT  13.505 0.850 13.860 1.080 ;
        RECT  13.505 2.880 13.800 3.220 ;
        RECT  13.340 0.850 13.505 3.220 ;
        RECT  13.275 0.850 13.340 3.165 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.405 4.465 2.075 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.150 1.235 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 -0.400 16.500 0.400 ;
        RECT  15.980 -0.400 16.320 0.575 ;
        RECT  15.000 -0.400 15.980 0.400 ;
        RECT  14.660 -0.400 15.000 0.575 ;
        RECT  13.400 -0.400 14.660 0.400 ;
        RECT  13.060 -0.400 13.400 0.575 ;
        RECT  11.440 -0.400 13.060 0.400 ;
        RECT  11.100 -0.400 11.440 1.270 ;
        RECT  8.825 -0.400 11.100 0.400 ;
        RECT  8.485 -0.400 8.825 1.440 ;
        RECT  6.660 -0.400 8.485 0.400 ;
        RECT  6.320 -0.400 6.660 1.270 ;
        RECT  3.140 -0.400 6.320 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.210 -0.400 2.800 0.400 ;
        RECT  1.210 1.440 1.240 1.780 ;
        RECT  0.870 -0.400 1.210 1.780 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.180 4.640 16.500 5.440 ;
        RECT  15.755 4.465 16.180 5.440 ;
        RECT  14.560 4.640 15.755 5.440 ;
        RECT  14.220 4.465 14.560 5.440 ;
        RECT  12.580 4.640 14.220 5.440 ;
        RECT  10.830 4.465 12.580 5.440 ;
        RECT  8.510 4.640 10.830 5.440 ;
        RECT  8.170 4.465 8.510 5.440 ;
        RECT  4.100 4.640 8.170 5.440 ;
        RECT  3.760 4.410 4.100 5.440 ;
        RECT  1.545 4.640 3.760 5.440 ;
        RECT  1.160 4.465 1.545 5.440 ;
        RECT  0.000 4.640 1.160 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.790 3.995 15.130 4.360 ;
        RECT  14.765 3.995 14.790 4.225 ;
        RECT  14.535 1.590 14.765 4.225 ;
        RECT  14.200 1.590 14.535 1.820 ;
        RECT  13.800 3.995 14.535 4.225 ;
        RECT  14.070 2.340 14.300 3.680 ;
        RECT  13.860 1.480 14.200 1.820 ;
        RECT  13.775 2.340 14.070 2.570 ;
        RECT  12.615 3.450 14.070 3.680 ;
        RECT  13.690 3.995 13.800 4.370 ;
        RECT  13.460 3.910 13.690 4.370 ;
        RECT  12.280 3.910 13.460 4.140 ;
        RECT  12.385 1.565 12.615 3.680 ;
        RECT  12.240 1.565 12.385 1.795 ;
        RECT  11.670 3.415 12.385 3.680 ;
        RECT  11.900 1.145 12.240 1.795 ;
        RECT  11.750 2.350 12.090 2.690 ;
        RECT  10.770 1.565 11.900 1.795 ;
        RECT  9.940 2.405 11.750 2.635 ;
        RECT  11.560 3.360 11.670 3.700 ;
        RECT  11.330 3.360 11.560 3.960 ;
        RECT  9.850 3.730 11.330 3.960 ;
        RECT  10.540 1.160 10.770 1.795 ;
        RECT  10.160 1.160 10.540 1.390 ;
        RECT  9.820 1.050 10.160 1.390 ;
        RECT  9.830 2.405 9.940 3.160 ;
        RECT  9.510 3.440 9.850 4.250 ;
        RECT  9.600 1.720 9.830 3.160 ;
        RECT  8.030 1.720 9.600 1.950 ;
        RECT  8.970 2.930 9.600 3.160 ;
        RECT  9.195 2.190 9.250 2.530 ;
        RECT  8.910 2.190 9.195 2.535 ;
        RECT  8.740 2.930 8.970 4.235 ;
        RECT  8.500 2.305 8.910 2.535 ;
        RECT  6.290 4.005 8.740 4.235 ;
        RECT  8.270 2.305 8.500 3.775 ;
        RECT  7.335 3.545 8.270 3.775 ;
        RECT  8.030 1.095 8.085 1.435 ;
        RECT  8.020 1.095 8.030 1.950 ;
        RECT  7.790 1.095 8.020 2.965 ;
        RECT  7.745 1.095 7.790 1.435 ;
        RECT  7.630 2.625 7.790 2.965 ;
        RECT  7.325 0.965 7.380 1.305 ;
        RECT  7.325 2.270 7.335 3.775 ;
        RECT  7.105 0.965 7.325 3.775 ;
        RECT  7.095 0.965 7.105 2.510 ;
        RECT  7.040 0.965 7.095 1.305 ;
        RECT  6.225 2.170 7.095 2.510 ;
        RECT  6.480 1.500 6.820 1.840 ;
        RECT  5.995 1.555 6.480 1.785 ;
        RECT  6.005 3.695 6.290 4.235 ;
        RECT  5.950 3.695 6.005 4.045 ;
        RECT  5.765 1.545 5.995 3.430 ;
        RECT  5.535 3.695 5.950 3.925 ;
        RECT  5.610 1.545 5.765 1.785 ;
        RECT  5.380 0.920 5.610 1.785 ;
        RECT  5.305 2.630 5.535 3.925 ;
        RECT  4.960 4.170 5.480 4.400 ;
        RECT  5.300 0.920 5.380 1.150 ;
        RECT  5.070 2.630 5.305 2.860 ;
        RECT  4.960 0.810 5.300 1.150 ;
        RECT  4.735 3.260 5.075 3.600 ;
        RECT  4.840 1.380 5.070 2.860 ;
        RECT  4.730 3.920 4.960 4.400 ;
        RECT  4.730 1.380 4.840 1.720 ;
        RECT  3.070 3.315 4.735 3.545 ;
        RECT  3.530 3.920 4.730 4.150 ;
        RECT  4.160 0.750 4.500 1.090 ;
        RECT  2.555 0.810 4.160 1.040 ;
        RECT  3.505 1.345 3.550 1.575 ;
        RECT  3.300 3.920 3.530 4.410 ;
        RECT  3.210 1.270 3.505 1.575 ;
        RECT  2.035 4.180 3.300 4.410 ;
        RECT  2.120 1.270 3.210 1.500 ;
        RECT  2.840 3.315 3.070 3.930 ;
        RECT  2.295 3.700 2.840 3.930 ;
        RECT  2.270 2.940 2.610 3.380 ;
        RECT  2.325 0.645 2.555 1.040 ;
        RECT  1.440 0.645 2.325 0.875 ;
        RECT  1.700 2.940 2.270 3.170 ;
        RECT  1.835 1.270 2.120 1.780 ;
        RECT  1.805 3.605 2.035 4.410 ;
        RECT  1.780 1.440 1.835 1.780 ;
        RECT  0.790 3.605 1.805 3.835 ;
        RECT  1.700 1.550 1.780 1.780 ;
        RECT  1.470 1.550 1.700 3.170 ;
        RECT  0.570 3.020 0.790 3.835 ;
        RECT  0.390 1.340 0.570 3.835 ;
        RECT  0.340 1.340 0.390 3.310 ;
        RECT  0.180 1.340 0.340 1.680 ;
    END
END SDFFNX2

MACRO SDFFNX1
    CLASS CORE ;
    FOREIGN SDFFNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.845 3.290 2.380 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.950 2.780 4.005 3.120 ;
        RECT  3.665 2.630 3.950 3.120 ;
        RECT  2.500 2.630 3.665 2.860 ;
        RECT  2.210 2.380 2.500 2.860 ;
        RECT  2.120 2.380 2.210 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.340 1.190 13.680 3.880 ;
        RECT  13.240 3.540 13.340 3.880 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 0.865 12.985 3.420 ;
        RECT  12.680 0.865 12.755 1.285 ;
        RECT  11.870 3.190 12.755 3.420 ;
        RECT  12.280 0.865 12.680 1.095 ;
        RECT  11.940 0.725 12.280 1.095 ;
        RECT  11.530 3.190 11.870 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 1.845 4.405 2.075 ;
        RECT  4.015 1.405 4.270 2.075 ;
        RECT  3.930 1.405 4.015 1.745 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.205 1.180 2.660 ;
        RECT  0.645 2.150 0.875 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.100 -0.400 13.860 0.400 ;
        RECT  12.760 -0.400 13.100 0.575 ;
        RECT  11.520 -0.400 12.760 0.400 ;
        RECT  11.180 -0.400 11.520 0.575 ;
        RECT  9.080 -0.400 11.180 0.400 ;
        RECT  8.740 -0.400 9.080 1.570 ;
        RECT  6.710 -0.400 8.740 0.400 ;
        RECT  6.370 -0.400 6.710 1.150 ;
        RECT  3.190 -0.400 6.370 0.400 ;
        RECT  2.850 -0.400 3.190 0.575 ;
        RECT  1.260 -0.400 2.850 0.400 ;
        RECT  1.260 1.345 1.530 1.685 ;
        RECT  1.190 -0.400 1.260 1.685 ;
        RECT  1.030 -0.400 1.190 1.630 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.820 4.640 13.860 5.440 ;
        RECT  12.480 4.410 12.820 5.440 ;
        RECT  11.110 4.640 12.480 5.440 ;
        RECT  10.770 4.465 11.110 5.440 ;
        RECT  8.435 4.640 10.770 5.440 ;
        RECT  8.095 4.465 8.435 5.440 ;
        RECT  4.035 4.640 8.095 5.440 ;
        RECT  3.695 4.410 4.035 5.440 ;
        RECT  0.735 4.640 3.695 5.440 ;
        RECT  0.395 4.410 0.735 5.440 ;
        RECT  0.000 4.640 0.395 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.365 2.005 12.510 2.430 ;
        RECT  12.135 1.470 12.365 2.955 ;
        RECT  11.980 1.470 12.135 1.810 ;
        RECT  10.990 2.725 12.135 2.955 ;
        RECT  11.555 2.040 11.895 2.380 ;
        RECT  11.760 4.030 11.870 4.370 ;
        RECT  11.530 3.970 11.760 4.370 ;
        RECT  11.520 2.040 11.555 2.270 ;
        RECT  10.990 3.970 11.530 4.200 ;
        RECT  11.290 1.440 11.520 2.270 ;
        RECT  10.190 1.440 11.290 1.835 ;
        RECT  10.760 2.180 10.990 4.200 ;
        RECT  10.650 2.180 10.760 2.520 ;
        RECT  9.580 0.670 10.740 0.900 ;
        RECT  9.960 1.440 10.190 4.230 ;
        RECT  9.850 4.000 9.960 4.230 ;
        RECT  9.510 4.000 9.850 4.340 ;
        RECT  9.505 2.820 9.730 3.160 ;
        RECT  9.505 0.670 9.580 2.070 ;
        RECT  9.350 0.670 9.505 3.615 ;
        RECT  9.275 1.840 9.350 3.615 ;
        RECT  8.250 1.840 9.275 2.070 ;
        RECT  8.910 3.385 9.275 3.615 ;
        RECT  8.775 2.380 9.005 3.135 ;
        RECT  8.680 3.385 8.910 4.235 ;
        RECT  8.440 2.905 8.775 3.135 ;
        RECT  6.230 4.005 8.680 4.235 ;
        RECT  8.210 2.905 8.440 3.775 ;
        RECT  7.970 1.120 8.250 2.070 ;
        RECT  7.400 3.545 8.210 3.775 ;
        RECT  7.910 1.120 7.970 3.130 ;
        RECT  7.740 1.840 7.910 3.130 ;
        RECT  7.630 2.790 7.740 3.130 ;
        RECT  7.455 0.810 7.510 1.150 ;
        RECT  7.400 0.810 7.455 2.400 ;
        RECT  7.225 0.810 7.400 3.775 ;
        RECT  7.170 0.810 7.225 1.150 ;
        RECT  7.130 2.060 7.225 3.775 ;
        RECT  6.220 2.060 7.130 2.400 ;
        RECT  6.655 1.385 6.995 1.725 ;
        RECT  5.935 1.440 6.655 1.670 ;
        RECT  6.120 3.950 6.230 4.290 ;
        RECT  5.890 3.720 6.120 4.290 ;
        RECT  5.705 0.805 5.935 3.490 ;
        RECT  5.475 3.720 5.890 3.950 ;
        RECT  5.010 0.805 5.705 1.035 ;
        RECT  5.015 4.180 5.535 4.410 ;
        RECT  5.245 2.820 5.475 3.950 ;
        RECT  5.015 2.820 5.245 3.050 ;
        RECT  5.015 1.390 5.070 1.730 ;
        RECT  4.785 1.390 5.015 3.050 ;
        RECT  4.675 3.320 5.015 3.660 ;
        RECT  4.785 3.920 5.015 4.410 ;
        RECT  4.730 1.390 4.785 1.730 ;
        RECT  3.455 3.920 4.785 4.150 ;
        RECT  2.990 3.375 4.675 3.605 ;
        RECT  4.210 0.750 4.550 1.090 ;
        RECT  2.605 0.810 4.210 1.040 ;
        RECT  2.380 1.345 3.595 1.575 ;
        RECT  3.225 3.920 3.455 4.410 ;
        RECT  1.895 4.180 3.225 4.410 ;
        RECT  2.760 3.375 2.990 3.930 ;
        RECT  2.145 3.700 2.760 3.930 ;
        RECT  2.375 0.645 2.605 1.040 ;
        RECT  1.890 3.095 2.530 3.325 ;
        RECT  2.270 1.345 2.380 1.770 ;
        RECT  1.490 0.645 2.375 0.875 ;
        RECT  2.095 1.345 2.270 2.150 ;
        RECT  2.040 1.430 2.095 2.150 ;
        RECT  1.890 1.920 2.040 2.150 ;
        RECT  1.665 3.605 1.895 4.410 ;
        RECT  1.660 1.920 1.890 3.325 ;
        RECT  0.570 3.605 1.665 3.835 ;
        RECT  1.520 2.885 1.660 3.325 ;
        RECT  0.410 1.430 0.750 1.770 ;
        RECT  0.380 3.020 0.570 3.835 ;
        RECT  0.380 1.540 0.410 1.770 ;
        RECT  0.150 1.540 0.380 3.835 ;
    END
END SDFFNX1

MACRO SDFFHQXL
    CLASS CORE ;
    FOREIGN SDFFHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.845 3.290 2.390 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 2.630 3.960 3.010 ;
        RECT  2.500 2.630 3.620 2.860 ;
        RECT  2.210 2.380 2.500 2.860 ;
        RECT  2.120 2.380 2.210 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.985 0.795 13.075 3.525 ;
        RECT  12.845 0.795 12.985 3.755 ;
        RECT  12.755 0.795 12.845 1.025 ;
        RECT  12.755 3.190 12.845 3.755 ;
        RECT  12.570 0.700 12.755 1.025 ;
        RECT  11.730 3.190 12.755 3.530 ;
        RECT  12.230 0.685 12.570 1.025 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 1.845 4.405 2.075 ;
        RECT  4.015 1.405 4.270 2.075 ;
        RECT  3.930 1.405 4.015 1.745 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.205 1.180 2.660 ;
        RECT  0.645 2.150 0.875 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.810 -0.400 13.200 0.400 ;
        RECT  11.470 -0.400 11.810 0.575 ;
        RECT  8.955 -0.400 11.470 0.400 ;
        RECT  8.725 -0.400 8.955 1.460 ;
        RECT  6.655 -0.400 8.725 0.400 ;
        RECT  6.425 -0.400 6.655 1.150 ;
        RECT  3.190 -0.400 6.425 0.400 ;
        RECT  2.850 -0.400 3.190 0.575 ;
        RECT  1.260 -0.400 2.850 0.400 ;
        RECT  1.260 1.290 1.580 1.630 ;
        RECT  1.240 -0.400 1.260 1.630 ;
        RECT  1.030 -0.400 1.240 1.520 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.270 4.640 13.200 5.440 ;
        RECT  10.930 4.465 11.270 5.440 ;
        RECT  8.435 4.640 10.930 5.440 ;
        RECT  8.095 4.465 8.435 5.440 ;
        RECT  4.340 4.640 8.095 5.440 ;
        RECT  4.000 4.410 4.340 5.440 ;
        RECT  1.100 4.640 4.000 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.565 1.460 12.610 1.800 ;
        RECT  12.335 1.460 12.565 2.960 ;
        RECT  12.270 1.460 12.335 1.800 ;
        RECT  11.280 2.730 12.335 2.960 ;
        RECT  11.810 2.040 12.105 2.380 ;
        RECT  11.690 4.005 12.030 4.400 ;
        RECT  11.580 1.605 11.810 2.380 ;
        RECT  11.280 4.005 11.690 4.235 ;
        RECT  10.595 1.605 11.580 1.835 ;
        RECT  11.050 2.180 11.280 4.235 ;
        RECT  10.940 2.180 11.050 2.520 ;
        RECT  9.415 0.875 11.030 1.105 ;
        RECT  10.365 1.370 10.595 4.240 ;
        RECT  10.050 4.010 10.365 4.240 ;
        RECT  9.905 1.335 10.135 3.670 ;
        RECT  9.710 4.010 10.050 4.350 ;
        RECT  9.645 1.335 9.905 1.675 ;
        RECT  9.275 3.440 9.905 3.670 ;
        RECT  9.445 1.905 9.675 3.190 ;
        RECT  9.415 1.905 9.445 2.135 ;
        RECT  8.775 2.960 9.445 3.190 ;
        RECT  9.185 0.875 9.415 2.135 ;
        RECT  9.045 3.440 9.275 4.185 ;
        RECT  8.545 1.905 9.185 2.135 ;
        RECT  8.720 2.380 9.060 2.720 ;
        RECT  8.545 2.960 8.775 4.235 ;
        RECT  8.315 2.490 8.720 2.720 ;
        RECT  8.315 1.765 8.545 2.135 ;
        RECT  6.240 4.005 8.545 4.235 ;
        RECT  8.200 1.765 8.315 1.995 ;
        RECT  8.085 2.490 8.315 3.775 ;
        RECT  8.005 1.170 8.210 1.510 ;
        RECT  7.265 3.545 8.085 3.775 ;
        RECT  7.915 0.630 8.005 1.510 ;
        RECT  7.855 0.630 7.915 1.615 ;
        RECT  7.775 0.630 7.855 3.130 ;
        RECT  7.685 1.225 7.775 3.130 ;
        RECT  7.625 1.385 7.685 3.130 ;
        RECT  7.265 0.810 7.455 1.155 ;
        RECT  7.225 0.810 7.265 3.775 ;
        RECT  7.035 0.925 7.225 3.775 ;
        RECT  6.560 2.240 7.035 2.470 ;
        RECT  6.575 1.455 6.805 1.800 ;
        RECT  5.935 1.455 6.575 1.685 ;
        RECT  6.220 2.130 6.560 2.470 ;
        RECT  6.230 3.920 6.240 4.235 ;
        RECT  5.890 3.920 6.230 4.290 ;
        RECT  5.705 0.805 5.935 3.680 ;
        RECT  5.475 3.920 5.890 4.150 ;
        RECT  5.010 0.805 5.705 1.035 ;
        RECT  5.245 2.820 5.475 4.150 ;
        RECT  5.070 2.820 5.245 3.050 ;
        RECT  3.770 3.920 5.245 4.150 ;
        RECT  4.840 1.390 5.070 3.050 ;
        RECT  4.675 3.320 5.015 3.660 ;
        RECT  4.730 1.390 4.840 1.730 ;
        RECT  3.310 3.430 4.675 3.660 ;
        RECT  4.210 0.750 4.550 1.090 ;
        RECT  2.605 0.810 4.210 1.040 ;
        RECT  3.540 3.920 3.770 4.410 ;
        RECT  2.380 1.355 3.595 1.585 ;
        RECT  1.895 4.180 3.540 4.410 ;
        RECT  3.080 3.430 3.310 3.930 ;
        RECT  2.145 3.700 3.080 3.930 ;
        RECT  1.890 3.095 2.850 3.325 ;
        RECT  2.375 0.645 2.605 1.040 ;
        RECT  2.270 1.355 2.380 1.750 ;
        RECT  1.490 0.645 2.375 0.875 ;
        RECT  2.040 1.355 2.270 2.145 ;
        RECT  1.890 1.915 2.040 2.145 ;
        RECT  1.665 3.605 1.895 4.410 ;
        RECT  1.660 1.915 1.890 3.325 ;
        RECT  0.570 3.605 1.665 3.835 ;
        RECT  1.520 2.885 1.660 3.225 ;
        RECT  0.410 1.410 0.750 1.750 ;
        RECT  0.380 3.020 0.570 3.835 ;
        RECT  0.380 1.520 0.410 1.750 ;
        RECT  0.150 1.520 0.380 3.835 ;
    END
END SDFFHQXL

MACRO SDFFHQX4
    CLASS CORE ;
    FOREIGN SDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFHQXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 1.820 3.320 2.240 ;
        RECT  2.860 1.820 3.200 2.295 ;
        RECT  2.780 1.820 2.860 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 2.490 3.870 2.830 ;
        RECT  2.630 2.525 3.530 2.755 ;
        RECT  2.400 2.380 2.630 2.755 ;
        RECT  2.010 2.380 2.400 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 1.820 16.360 3.220 ;
        RECT  15.990 1.365 16.330 3.220 ;
        RECT  15.980 1.820 15.990 3.220 ;
        RECT  15.750 2.820 15.980 3.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 1.495 4.410 1.845 ;
        RECT  4.385 2.405 4.405 2.635 ;
        RECT  4.150 1.495 4.385 2.635 ;
        RECT  4.070 1.495 4.150 1.835 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 2.200 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.970 -0.400 17.160 0.400 ;
        RECT  16.630 -0.400 16.970 0.965 ;
        RECT  15.690 -0.400 16.630 0.400 ;
        RECT  15.350 -0.400 15.690 0.955 ;
        RECT  14.190 -0.400 15.350 0.400 ;
        RECT  13.850 -0.400 14.190 0.575 ;
        RECT  12.375 -0.400 13.850 0.400 ;
        RECT  12.145 -0.400 12.375 1.270 ;
        RECT  9.235 -0.400 12.145 0.400 ;
        RECT  9.005 -0.400 9.235 1.370 ;
        RECT  6.740 -0.400 9.005 0.400 ;
        RECT  6.400 -0.400 6.740 1.270 ;
        RECT  3.220 -0.400 6.400 0.400 ;
        RECT  2.880 -0.400 3.220 0.575 ;
        RECT  1.290 -0.400 2.880 0.400 ;
        RECT  1.290 1.445 1.320 1.785 ;
        RECT  0.950 -0.400 1.290 1.785 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.735 4.640 17.160 5.440 ;
        RECT  16.395 4.090 16.735 5.440 ;
        RECT  15.405 4.640 16.395 5.440 ;
        RECT  15.065 4.465 15.405 5.440 ;
        RECT  14.060 4.640 15.065 5.440 ;
        RECT  11.670 4.465 14.060 5.440 ;
        RECT  9.050 4.640 11.670 5.440 ;
        RECT  8.710 4.465 9.050 5.440 ;
        RECT  5.640 4.640 8.710 5.440 ;
        RECT  5.300 4.465 5.640 5.440 ;
        RECT  1.285 4.640 5.300 5.440 ;
        RECT  0.945 4.465 1.285 5.440 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.960 1.110 14.990 1.450 ;
        RECT  14.730 1.110 14.960 3.810 ;
        RECT  14.650 1.110 14.730 2.400 ;
        RECT  14.485 3.470 14.730 3.810 ;
        RECT  14.105 2.060 14.650 2.400 ;
        RECT  13.865 2.730 14.500 3.070 ;
        RECT  13.635 1.500 13.865 3.720 ;
        RECT  13.230 1.500 13.635 1.730 ;
        RECT  12.825 3.490 13.635 3.720 ;
        RECT  13.020 1.960 13.250 3.225 ;
        RECT  12.890 0.630 13.230 1.730 ;
        RECT  11.450 1.960 13.020 2.190 ;
        RECT  12.360 2.995 13.020 3.225 ;
        RECT  11.915 1.500 12.890 1.730 ;
        RECT  12.595 3.490 12.825 4.235 ;
        RECT  12.450 2.425 12.790 2.765 ;
        RECT  10.530 4.005 12.595 4.235 ;
        RECT  11.900 2.535 12.450 2.765 ;
        RECT  12.130 2.995 12.360 3.770 ;
        RECT  9.810 3.540 12.130 3.770 ;
        RECT  11.685 0.935 11.915 1.730 ;
        RECT  11.670 2.535 11.900 3.305 ;
        RECT  10.730 0.935 11.685 1.165 ;
        RECT  10.240 3.075 11.670 3.305 ;
        RECT  11.220 1.460 11.450 2.190 ;
        RECT  11.100 2.505 11.440 2.845 ;
        RECT  11.110 1.460 11.220 1.800 ;
        RECT  10.020 1.570 11.110 1.800 ;
        RECT  10.705 2.510 11.100 2.740 ;
        RECT  10.390 0.935 10.730 1.275 ;
        RECT  10.475 2.060 10.705 2.740 ;
        RECT  10.190 4.005 10.530 4.345 ;
        RECT  9.570 2.060 10.475 2.290 ;
        RECT  9.900 2.540 10.240 3.305 ;
        RECT  9.790 1.030 10.020 1.800 ;
        RECT  8.950 3.075 9.900 3.305 ;
        RECT  9.470 3.540 9.810 3.880 ;
        RECT  9.670 1.030 9.790 1.370 ;
        RECT  9.460 2.060 9.570 2.400 ;
        RECT  9.230 1.600 9.460 2.400 ;
        RECT  8.775 1.600 9.230 1.830 ;
        RECT  8.810 2.225 8.950 4.170 ;
        RECT  8.720 2.115 8.810 4.170 ;
        RECT  8.545 0.665 8.775 1.830 ;
        RECT  8.470 2.115 8.720 2.455 ;
        RECT  6.230 3.940 8.720 4.170 ;
        RECT  7.460 0.665 8.545 0.895 ;
        RECT  8.380 3.315 8.490 3.655 ;
        RECT  8.240 2.850 8.380 3.655 ;
        RECT  8.240 1.130 8.315 1.690 ;
        RECT  8.150 1.130 8.240 3.655 ;
        RECT  8.085 1.130 8.150 3.080 ;
        RECT  8.010 1.460 8.085 3.080 ;
        RECT  7.665 1.905 8.010 2.245 ;
        RECT  7.445 3.320 7.785 3.660 ;
        RECT  7.435 0.665 7.460 1.485 ;
        RECT  7.435 3.320 7.445 3.605 ;
        RECT  7.230 0.665 7.435 3.605 ;
        RECT  7.205 1.145 7.230 3.605 ;
        RECT  7.120 1.145 7.205 1.485 ;
        RECT  6.440 2.570 7.205 2.910 ;
        RECT  6.635 1.890 6.975 2.230 ;
        RECT  5.810 1.890 6.635 2.120 ;
        RECT  5.890 3.940 6.230 4.280 ;
        RECT  5.350 3.945 5.890 4.175 ;
        RECT  5.580 0.685 5.810 3.590 ;
        RECT  5.040 0.685 5.580 0.915 ;
        RECT  5.120 1.500 5.350 4.175 ;
        RECT  5.100 1.500 5.120 1.730 ;
        RECT  4.365 3.945 5.120 4.175 ;
        RECT  4.760 1.390 5.100 1.730 ;
        RECT  4.550 3.260 4.890 3.600 ;
        RECT  4.240 0.670 4.580 1.035 ;
        RECT  3.860 3.370 4.550 3.600 ;
        RECT  4.135 3.945 4.365 4.410 ;
        RECT  1.870 0.805 4.240 1.035 ;
        RECT  1.840 4.180 4.135 4.410 ;
        RECT  3.630 3.370 3.860 3.930 ;
        RECT  2.210 1.335 3.630 1.565 ;
        RECT  2.070 3.700 3.630 3.930 ;
        RECT  2.310 3.040 2.650 3.380 ;
        RECT  1.940 3.040 2.310 3.270 ;
        RECT  2.100 1.335 2.210 1.785 ;
        RECT  1.870 1.335 2.100 2.150 ;
        RECT  1.780 2.905 1.940 3.270 ;
        RECT  1.520 0.645 1.870 1.035 ;
        RECT  1.780 1.920 1.870 2.150 ;
        RECT  1.610 3.685 1.840 4.410 ;
        RECT  1.550 1.920 1.780 3.270 ;
        RECT  0.520 3.685 1.610 3.915 ;
        RECT  0.350 1.445 0.600 1.785 ;
        RECT  0.465 3.105 0.520 3.915 ;
        RECT  0.350 2.890 0.465 3.915 ;
        RECT  0.260 1.445 0.350 3.915 ;
        RECT  0.180 1.550 0.260 3.915 ;
        RECT  0.120 1.550 0.180 3.120 ;
    END
END SDFFHQX4

MACRO SDFFHQX2
    CLASS CORE ;
    FOREIGN SDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFHQXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.980 1.820 3.160 2.100 ;
        RECT  2.470 1.730 2.980 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.995 2.720 4.105 3.060 ;
        RECT  3.765 2.410 3.995 3.060 ;
        RECT  2.500 2.410 3.765 2.640 ;
        RECT  2.120 2.380 2.500 2.665 ;
        RECT  2.050 2.385 2.120 2.665 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.540 0.700 14.880 1.040 ;
        RECT  14.165 0.810 14.540 1.040 ;
        RECT  14.165 2.940 14.380 3.220 ;
        RECT  13.935 0.810 14.165 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.405 4.465 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.150 1.235 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.640 -0.400 15.840 0.400 ;
        RECT  15.300 -0.400 15.640 0.950 ;
        RECT  14.080 -0.400 15.300 0.400 ;
        RECT  13.740 -0.400 14.080 0.575 ;
        RECT  12.065 -0.400 13.740 0.400 ;
        RECT  11.835 -0.400 12.065 1.075 ;
        RECT  8.960 -0.400 11.835 0.400 ;
        RECT  8.620 -0.400 8.960 1.355 ;
        RECT  6.660 -0.400 8.620 0.400 ;
        RECT  6.320 -0.400 6.660 1.270 ;
        RECT  3.140 -0.400 6.320 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.210 -0.400 2.800 0.400 ;
        RECT  1.210 1.440 1.240 1.780 ;
        RECT  0.870 -0.400 1.210 1.780 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.980 4.640 15.840 5.440 ;
        RECT  14.640 4.465 14.980 5.440 ;
        RECT  13.000 4.640 14.640 5.440 ;
        RECT  11.250 4.465 13.000 5.440 ;
        RECT  8.570 4.640 11.250 5.440 ;
        RECT  8.230 4.465 8.570 5.440 ;
        RECT  4.100 4.640 8.230 5.440 ;
        RECT  3.760 4.410 4.100 5.440 ;
        RECT  1.520 4.640 3.760 5.440 ;
        RECT  1.180 4.465 1.520 5.440 ;
        RECT  0.000 4.640 1.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.075 1.570 15.305 4.140 ;
        RECT  14.880 1.570 15.075 1.800 ;
        RECT  14.220 3.910 15.075 4.140 ;
        RECT  14.540 1.460 14.880 1.800 ;
        RECT  14.610 2.285 14.840 3.680 ;
        RECT  13.705 3.450 14.610 3.680 ;
        RECT  13.875 3.910 14.220 4.370 ;
        RECT  13.040 3.910 13.875 4.140 ;
        RECT  13.475 1.500 13.705 3.680 ;
        RECT  12.920 1.500 13.475 1.730 ;
        RECT  12.090 3.360 13.475 3.590 ;
        RECT  13.015 1.960 13.245 3.130 ;
        RECT  12.700 3.850 13.040 4.190 ;
        RECT  11.105 1.960 13.015 2.190 ;
        RECT  10.830 2.900 13.015 3.130 ;
        RECT  12.580 1.165 12.920 1.730 ;
        RECT  10.110 2.420 12.710 2.650 ;
        RECT  11.565 1.500 12.580 1.730 ;
        RECT  11.980 3.360 12.090 3.700 ;
        RECT  11.750 3.360 11.980 4.190 ;
        RECT  10.110 3.960 11.750 4.190 ;
        RECT  11.335 0.640 11.565 1.730 ;
        RECT  10.445 0.640 11.335 0.870 ;
        RECT  10.875 1.100 11.105 2.190 ;
        RECT  9.720 1.445 10.875 1.675 ;
        RECT  10.600 2.900 10.830 3.730 ;
        RECT  10.490 3.390 10.600 3.730 ;
        RECT  9.335 3.390 10.490 3.620 ;
        RECT  10.215 0.640 10.445 1.215 ;
        RECT  10.100 0.985 10.215 1.215 ;
        RECT  10.000 2.420 10.110 3.160 ;
        RECT  9.770 3.850 10.110 4.190 ;
        RECT  9.770 1.905 10.000 3.160 ;
        RECT  8.150 1.905 9.770 2.135 ;
        RECT  8.875 2.930 9.770 3.160 ;
        RECT  9.490 1.100 9.720 1.675 ;
        RECT  9.380 1.100 9.490 1.440 ;
        RECT  9.105 3.390 9.335 3.730 ;
        RECT  8.415 2.365 9.250 2.595 ;
        RECT  8.645 2.930 8.875 4.235 ;
        RECT  6.330 4.005 8.645 4.235 ;
        RECT  8.185 2.365 8.415 3.775 ;
        RECT  7.405 3.545 8.185 3.775 ;
        RECT  8.015 1.105 8.160 1.445 ;
        RECT  7.920 0.630 8.015 1.445 ;
        RECT  7.920 2.365 7.955 2.965 ;
        RECT  7.725 0.630 7.920 2.965 ;
        RECT  7.690 0.630 7.725 2.595 ;
        RECT  7.655 0.630 7.690 0.860 ;
        RECT  7.175 0.950 7.405 3.775 ;
        RECT  6.265 2.160 7.175 2.500 ;
        RECT  6.035 1.545 6.820 1.775 ;
        RECT  6.325 3.920 6.330 4.280 ;
        RECT  5.990 3.890 6.325 4.280 ;
        RECT  5.805 1.545 6.035 3.600 ;
        RECT  5.575 3.890 5.990 4.150 ;
        RECT  5.610 1.545 5.805 1.775 ;
        RECT  5.380 0.920 5.610 1.775 ;
        RECT  5.345 2.600 5.575 4.150 ;
        RECT  5.300 0.920 5.380 1.150 ;
        RECT  5.065 2.600 5.345 2.830 ;
        RECT  3.530 3.920 5.345 4.150 ;
        RECT  4.960 0.810 5.300 1.150 ;
        RECT  4.775 3.230 5.115 3.570 ;
        RECT  5.065 1.380 5.070 1.720 ;
        RECT  4.835 1.380 5.065 2.830 ;
        RECT  4.730 1.380 4.835 1.720 ;
        RECT  3.070 3.340 4.775 3.570 ;
        RECT  4.160 0.750 4.500 1.090 ;
        RECT  2.555 0.810 4.160 1.040 ;
        RECT  3.210 1.270 3.550 1.565 ;
        RECT  3.300 3.920 3.530 4.410 ;
        RECT  1.980 4.180 3.300 4.410 ;
        RECT  2.120 1.270 3.210 1.500 ;
        RECT  2.840 3.340 3.070 3.930 ;
        RECT  2.295 3.700 2.840 3.930 ;
        RECT  2.270 3.040 2.610 3.380 ;
        RECT  2.325 0.645 2.555 1.040 ;
        RECT  1.440 0.645 2.325 0.875 ;
        RECT  2.080 3.040 2.270 3.270 ;
        RECT  1.835 1.270 2.120 1.780 ;
        RECT  1.700 2.940 2.080 3.270 ;
        RECT  1.750 3.605 1.980 4.410 ;
        RECT  1.780 1.440 1.835 1.780 ;
        RECT  1.700 1.550 1.780 1.780 ;
        RECT  0.790 3.605 1.750 3.835 ;
        RECT  1.580 1.550 1.700 3.270 ;
        RECT  1.470 1.550 1.580 3.170 ;
        RECT  0.570 3.020 0.790 3.835 ;
        RECT  0.390 1.340 0.570 3.835 ;
        RECT  0.340 1.340 0.390 3.310 ;
        RECT  0.180 1.340 0.340 1.680 ;
    END
END SDFFHQX2

MACRO SDFFHQX1
    CLASS CORE ;
    FOREIGN SDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFHQXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.820 3.485 2.300 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 2.580 3.960 3.120 ;
        RECT  2.500 2.580 3.620 2.810 ;
        RECT  2.125 2.380 2.500 2.810 ;
        RECT  2.120 2.380 2.125 2.660 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.985 0.790 13.075 3.525 ;
        RECT  12.845 0.790 12.985 3.755 ;
        RECT  12.755 0.790 12.845 1.020 ;
        RECT  12.755 3.190 12.845 3.755 ;
        RECT  12.570 0.700 12.755 1.020 ;
        RECT  11.690 3.190 12.755 3.530 ;
        RECT  12.230 0.680 12.570 1.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 1.845 4.405 2.075 ;
        RECT  4.015 1.405 4.270 2.075 ;
        RECT  3.930 1.405 4.015 1.745 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.205 1.180 2.660 ;
        RECT  0.645 2.150 0.875 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.810 -0.400 13.200 0.400 ;
        RECT  11.470 -0.400 11.810 0.575 ;
        RECT  8.955 -0.400 11.470 0.400 ;
        RECT  8.725 -0.400 8.955 1.460 ;
        RECT  6.710 -0.400 8.725 0.400 ;
        RECT  6.370 -0.400 6.710 1.150 ;
        RECT  3.190 -0.400 6.370 0.400 ;
        RECT  2.850 -0.400 3.190 0.575 ;
        RECT  1.260 -0.400 2.850 0.400 ;
        RECT  1.260 1.290 1.530 1.630 ;
        RECT  1.190 -0.400 1.260 1.630 ;
        RECT  1.030 -0.400 1.190 1.520 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.790 4.640 13.200 5.440 ;
        RECT  12.450 4.410 12.790 5.440 ;
        RECT  11.270 4.640 12.450 5.440 ;
        RECT  10.930 4.465 11.270 5.440 ;
        RECT  8.340 4.640 10.930 5.440 ;
        RECT  7.060 4.465 8.340 5.440 ;
        RECT  4.340 4.640 7.060 5.440 ;
        RECT  4.000 4.410 4.340 5.440 ;
        RECT  1.100 4.640 4.000 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.380 1.460 12.610 2.960 ;
        RECT  12.270 1.460 12.380 1.800 ;
        RECT  11.280 2.730 12.380 2.960 ;
        RECT  11.875 2.040 12.105 2.380 ;
        RECT  11.730 4.115 12.030 4.345 ;
        RECT  11.810 2.040 11.875 2.270 ;
        RECT  11.580 1.605 11.810 2.270 ;
        RECT  11.500 4.005 11.730 4.345 ;
        RECT  10.595 1.605 11.580 1.835 ;
        RECT  11.280 4.005 11.500 4.235 ;
        RECT  11.050 2.180 11.280 4.235 ;
        RECT  10.940 2.180 11.050 2.520 ;
        RECT  10.690 0.820 11.030 1.160 ;
        RECT  9.415 0.875 10.690 1.105 ;
        RECT  10.365 1.440 10.595 4.235 ;
        RECT  10.010 4.005 10.365 4.235 ;
        RECT  9.905 1.445 10.135 3.710 ;
        RECT  9.670 4.005 10.010 4.345 ;
        RECT  9.875 1.445 9.905 1.675 ;
        RECT  9.235 3.480 9.905 3.710 ;
        RECT  9.645 1.335 9.875 1.675 ;
        RECT  9.505 2.820 9.675 3.235 ;
        RECT  9.415 1.910 9.505 3.235 ;
        RECT  9.275 0.875 9.415 3.235 ;
        RECT  9.185 0.875 9.275 2.140 ;
        RECT  8.775 3.005 9.275 3.235 ;
        RECT  9.005 3.480 9.235 4.185 ;
        RECT  8.200 1.765 9.185 1.995 ;
        RECT  8.315 2.380 9.005 2.735 ;
        RECT  8.545 3.005 8.775 4.235 ;
        RECT  6.230 4.005 8.545 4.235 ;
        RECT  8.085 2.380 8.315 3.775 ;
        RECT  8.060 1.170 8.210 1.510 ;
        RECT  7.320 3.545 8.085 3.775 ;
        RECT  7.950 0.630 8.060 1.510 ;
        RECT  7.855 0.630 7.950 1.615 ;
        RECT  7.720 0.630 7.855 3.130 ;
        RECT  7.625 1.385 7.720 3.130 ;
        RECT  7.320 0.810 7.455 1.155 ;
        RECT  7.225 0.810 7.320 3.775 ;
        RECT  7.090 0.925 7.225 3.775 ;
        RECT  6.450 2.130 7.090 2.470 ;
        RECT  6.520 1.460 6.860 1.800 ;
        RECT  5.935 1.570 6.520 1.800 ;
        RECT  5.890 3.950 6.230 4.290 ;
        RECT  5.705 0.805 5.935 3.680 ;
        RECT  5.475 3.950 5.890 4.180 ;
        RECT  5.350 0.805 5.705 1.090 ;
        RECT  5.245 1.500 5.475 4.180 ;
        RECT  5.010 0.750 5.350 1.090 ;
        RECT  5.070 1.500 5.245 1.730 ;
        RECT  3.770 3.950 5.245 4.180 ;
        RECT  4.730 1.390 5.070 1.730 ;
        RECT  4.675 3.320 5.015 3.660 ;
        RECT  3.310 3.430 4.675 3.660 ;
        RECT  4.210 0.750 4.550 1.090 ;
        RECT  2.605 0.860 4.210 1.090 ;
        RECT  3.540 3.950 3.770 4.410 ;
        RECT  2.380 1.345 3.595 1.575 ;
        RECT  1.895 4.180 3.540 4.410 ;
        RECT  3.080 3.430 3.310 3.930 ;
        RECT  2.145 3.700 3.080 3.930 ;
        RECT  2.390 3.040 2.730 3.380 ;
        RECT  2.375 0.645 2.605 1.090 ;
        RECT  1.890 3.040 2.390 3.270 ;
        RECT  2.040 1.345 2.380 1.770 ;
        RECT  1.490 0.645 2.375 0.875 ;
        RECT  1.990 1.540 2.040 1.770 ;
        RECT  1.890 1.540 1.990 2.145 ;
        RECT  1.665 3.605 1.895 4.410 ;
        RECT  1.760 1.540 1.890 3.270 ;
        RECT  1.660 1.915 1.760 3.270 ;
        RECT  0.570 3.605 1.665 3.835 ;
        RECT  1.520 2.885 1.660 3.270 ;
        RECT  0.410 1.430 0.750 1.770 ;
        RECT  0.380 3.020 0.570 3.835 ;
        RECT  0.380 1.540 0.410 1.770 ;
        RECT  0.150 1.540 0.380 3.835 ;
    END
END SDFFHQX1

MACRO SDFFXL
    CLASS CORE ;
    FOREIGN SDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 1.820 3.160 2.100 ;
        RECT  2.365 1.730 2.695 2.100 ;
        RECT  2.310 1.730 2.365 1.960 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.570 2.600 3.910 2.940 ;
        RECT  3.180 2.600 3.570 2.830 ;
        RECT  2.950 2.380 3.180 2.830 ;
        RECT  2.215 2.380 2.950 2.660 ;
        RECT  1.875 2.345 2.215 2.685 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.985 3.515 13.020 3.855 ;
        RECT  12.820 1.185 12.985 3.855 ;
        RECT  12.755 1.090 12.820 3.855 ;
        RECT  12.480 1.090 12.755 1.430 ;
        RECT  12.680 3.515 12.755 3.855 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.975 0.685 11.980 1.040 ;
        RECT  11.635 0.630 11.975 1.040 ;
        RECT  11.655 2.155 11.840 3.440 ;
        RECT  11.610 2.155 11.655 3.550 ;
        RECT  11.395 0.810 11.635 1.040 ;
        RECT  11.395 2.155 11.610 2.385 ;
        RECT  11.315 3.210 11.610 3.550 ;
        RECT  11.165 0.810 11.395 2.385 ;
        RECT  10.775 1.260 11.165 1.540 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.810 1.320 4.150 2.075 ;
        RECT  3.515 1.845 3.810 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.255 1.180 2.660 ;
        RECT  0.800 2.200 0.875 2.660 ;
        RECT  0.645 2.200 0.800 2.655 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.780 -0.400 13.200 0.400 ;
        RECT  12.440 -0.400 12.780 0.575 ;
        RECT  11.215 -0.400 12.440 0.400 ;
        RECT  10.875 -0.400 11.215 0.575 ;
        RECT  8.775 -0.400 10.875 0.400 ;
        RECT  8.435 -0.400 8.775 1.510 ;
        RECT  6.470 -0.400 8.435 0.400 ;
        RECT  6.130 -0.400 6.470 1.150 ;
        RECT  3.070 -0.400 6.130 0.400 ;
        RECT  2.730 -0.400 3.070 0.575 ;
        RECT  1.140 -0.400 2.730 0.400 ;
        RECT  1.140 1.290 1.320 1.630 ;
        RECT  0.980 -0.400 1.140 1.630 ;
        RECT  0.910 -0.400 0.980 1.575 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.315 4.640 13.200 5.440 ;
        RECT  11.975 4.410 12.315 5.440 ;
        RECT  10.850 4.640 11.975 5.440 ;
        RECT  10.510 4.465 10.850 5.440 ;
        RECT  8.365 4.640 10.510 5.440 ;
        RECT  7.085 4.465 8.365 5.440 ;
        RECT  4.020 4.640 7.085 5.440 ;
        RECT  3.680 4.410 4.020 5.440 ;
        RECT  1.100 4.640 3.680 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.220 1.685 12.450 4.180 ;
        RECT  11.960 1.685 12.220 1.915 ;
        RECT  11.735 3.950 12.220 4.180 ;
        RECT  11.730 1.360 11.960 1.915 ;
        RECT  11.505 3.950 11.735 4.350 ;
        RECT  11.240 4.005 11.505 4.350 ;
        RECT  11.035 2.615 11.375 2.955 ;
        RECT  10.420 4.005 11.240 4.235 ;
        RECT  10.880 2.615 11.035 2.845 ;
        RECT  10.650 1.840 10.880 2.845 ;
        RECT  10.055 1.840 10.650 2.070 ;
        RECT  10.190 2.505 10.420 4.235 ;
        RECT  9.295 0.670 10.335 0.900 ;
        RECT  9.945 1.270 10.055 2.070 ;
        RECT  9.715 1.270 9.945 4.150 ;
        RECT  9.685 3.920 9.715 4.150 ;
        RECT  9.345 3.920 9.685 4.260 ;
        RECT  9.295 2.920 9.315 3.260 ;
        RECT  9.205 0.670 9.295 3.260 ;
        RECT  9.115 0.670 9.205 3.595 ;
        RECT  9.065 0.670 9.115 4.235 ;
        RECT  8.135 1.740 9.065 1.970 ;
        RECT  8.975 2.920 9.065 4.235 ;
        RECT  8.885 3.365 8.975 4.235 ;
        RECT  6.195 4.005 8.885 4.235 ;
        RECT  8.605 2.200 8.830 2.545 ;
        RECT  8.440 2.200 8.605 3.135 ;
        RECT  8.375 2.200 8.440 3.775 ;
        RECT  8.210 2.905 8.375 3.775 ;
        RECT  6.920 3.545 8.210 3.775 ;
        RECT  7.905 1.740 8.135 2.510 ;
        RECT  7.875 1.170 7.975 1.510 ;
        RECT  7.675 0.630 7.875 1.510 ;
        RECT  7.675 2.780 7.770 3.120 ;
        RECT  7.445 0.630 7.675 3.120 ;
        RECT  7.430 2.780 7.445 3.120 ;
        RECT  6.985 0.810 7.215 2.425 ;
        RECT  6.920 2.195 6.985 2.425 ;
        RECT  6.690 2.195 6.920 3.775 ;
        RECT  6.410 1.590 6.750 1.930 ;
        RECT  6.310 2.400 6.690 2.740 ;
        RECT  5.890 1.590 6.410 1.820 ;
        RECT  5.855 3.950 6.195 4.290 ;
        RECT  5.795 0.850 5.890 1.820 ;
        RECT  5.335 3.950 5.855 4.180 ;
        RECT  5.565 0.850 5.795 3.680 ;
        RECT  5.110 0.850 5.565 1.080 ;
        RECT  5.105 2.820 5.335 4.180 ;
        RECT  4.770 0.740 5.110 1.080 ;
        RECT  4.765 2.820 5.105 3.050 ;
        RECT  3.450 3.950 5.105 4.180 ;
        RECT  4.535 3.320 4.875 3.660 ;
        RECT  4.535 1.390 4.765 3.050 ;
        RECT  2.990 3.375 4.535 3.605 ;
        RECT  4.050 0.750 4.390 1.090 ;
        RECT  2.485 0.810 4.050 1.040 ;
        RECT  3.220 3.950 3.450 4.410 ;
        RECT  2.960 1.270 3.350 1.575 ;
        RECT  1.730 4.180 3.220 4.410 ;
        RECT  2.760 3.375 2.990 3.930 ;
        RECT  2.065 1.270 2.960 1.500 ;
        RECT  2.095 3.700 2.760 3.930 ;
        RECT  2.255 0.645 2.485 1.040 ;
        RECT  2.135 3.050 2.475 3.450 ;
        RECT  1.370 0.645 2.255 0.875 ;
        RECT  1.860 3.050 2.135 3.280 ;
        RECT  1.835 1.270 2.065 2.095 ;
        RECT  1.645 2.940 1.860 3.280 ;
        RECT  1.645 1.865 1.835 2.095 ;
        RECT  1.500 3.935 1.730 4.410 ;
        RECT  1.415 1.865 1.645 3.280 ;
        RECT  0.540 3.935 1.500 4.165 ;
        RECT  0.380 3.015 0.540 4.165 ;
        RECT  0.380 1.430 0.520 1.770 ;
        RECT  0.310 1.430 0.380 4.165 ;
        RECT  0.150 1.430 0.310 3.360 ;
    END
END SDFFXL

MACRO SDFFX4
    CLASS CORE ;
    FOREIGN SDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 1.820 3.320 2.240 ;
        RECT  2.860 1.820 3.200 2.295 ;
        RECT  2.780 1.820 2.860 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 2.490 3.870 2.830 ;
        RECT  2.630 2.600 3.530 2.830 ;
        RECT  2.400 2.380 2.630 2.830 ;
        RECT  2.350 2.380 2.400 2.660 ;
        RECT  2.010 2.305 2.350 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.060 0.680 18.170 1.490 ;
        RECT  17.830 0.680 18.060 2.005 ;
        RECT  17.690 2.865 18.030 3.675 ;
        RECT  17.685 1.775 17.830 2.005 ;
        RECT  17.680 2.865 17.690 3.220 ;
        RECT  17.680 1.775 17.685 2.635 ;
        RECT  17.455 1.775 17.680 3.220 ;
        RECT  17.300 1.820 17.455 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.530 0.835 16.650 1.645 ;
        RECT  16.300 0.835 16.530 3.675 ;
        RECT  16.170 1.820 16.300 3.675 ;
        RECT  15.980 1.820 16.170 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.405 4.405 2.635 ;
        RECT  4.380 1.550 4.385 2.635 ;
        RECT  4.150 1.495 4.380 2.635 ;
        RECT  4.040 1.495 4.150 1.835 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 2.200 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.950 -0.400 19.140 0.400 ;
        RECT  18.610 -0.400 18.950 1.595 ;
        RECT  17.410 -0.400 18.610 0.400 ;
        RECT  17.070 -0.400 17.410 1.200 ;
        RECT  15.930 -0.400 17.070 0.400 ;
        RECT  15.590 -0.400 15.930 1.350 ;
        RECT  14.435 -0.400 15.590 0.400 ;
        RECT  14.205 -0.400 14.435 1.310 ;
        RECT  11.850 -0.400 14.205 0.400 ;
        RECT  11.510 -0.400 11.850 1.305 ;
        RECT  9.235 -0.400 11.510 0.400 ;
        RECT  9.005 -0.400 9.235 1.370 ;
        RECT  6.740 -0.400 9.005 0.400 ;
        RECT  6.400 -0.400 6.740 1.270 ;
        RECT  3.220 -0.400 6.400 0.400 ;
        RECT  2.880 -0.400 3.220 0.575 ;
        RECT  1.290 -0.400 2.880 0.400 ;
        RECT  1.290 1.445 1.320 1.785 ;
        RECT  0.980 -0.400 1.290 1.785 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.790 4.640 19.140 5.440 ;
        RECT  18.450 4.465 18.790 5.440 ;
        RECT  17.270 4.640 18.450 5.440 ;
        RECT  16.930 4.465 17.270 5.440 ;
        RECT  15.750 4.640 16.930 5.440 ;
        RECT  15.410 4.465 15.750 5.440 ;
        RECT  14.430 4.640 15.410 5.440 ;
        RECT  14.090 4.465 14.430 5.440 ;
        RECT  11.985 4.640 14.090 5.440 ;
        RECT  11.645 4.005 11.985 5.440 ;
        RECT  9.160 4.640 11.645 5.440 ;
        RECT  8.820 4.465 9.160 5.440 ;
        RECT  5.760 4.640 8.820 5.440 ;
        RECT  5.215 4.465 5.760 5.440 ;
        RECT  1.380 4.640 5.215 5.440 ;
        RECT  1.040 4.465 1.380 5.440 ;
        RECT  0.000 4.640 1.040 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.260 2.235 18.490 4.160 ;
        RECT  18.070 2.235 18.260 2.575 ;
        RECT  15.340 3.930 18.260 4.160 ;
        RECT  15.210 2.115 15.340 4.160 ;
        RECT  15.110 1.040 15.210 4.160 ;
        RECT  14.870 1.040 15.110 2.400 ;
        RECT  14.850 3.470 15.110 3.810 ;
        RECT  14.240 2.060 14.870 2.400 ;
        RECT  13.965 2.730 14.870 3.070 ;
        RECT  13.735 0.970 13.965 3.490 ;
        RECT  13.130 0.970 13.735 1.250 ;
        RECT  13.270 3.260 13.735 3.490 ;
        RECT  12.900 1.550 13.500 1.780 ;
        RECT  12.930 3.260 13.270 4.070 ;
        RECT  12.790 0.965 13.130 1.305 ;
        RECT  10.700 3.450 12.930 3.680 ;
        RECT  12.670 1.550 12.900 3.000 ;
        RECT  12.440 1.075 12.790 1.305 ;
        RECT  12.560 2.595 12.670 3.000 ;
        RECT  10.940 2.770 12.560 3.000 ;
        RECT  12.210 1.075 12.440 1.805 ;
        RECT  10.570 1.575 12.210 1.805 ;
        RECT  11.585 2.035 11.925 2.420 ;
        RECT  9.660 2.035 11.585 2.265 ;
        RECT  10.600 2.595 10.940 3.000 ;
        RECT  10.360 3.450 10.700 4.260 ;
        RECT  9.435 2.760 10.600 3.000 ;
        RECT  10.230 0.965 10.570 1.805 ;
        RECT  9.550 2.035 9.660 2.400 ;
        RECT  9.320 1.600 9.550 2.400 ;
        RECT  9.205 2.760 9.435 4.225 ;
        RECT  8.775 1.600 9.320 1.830 ;
        RECT  9.085 2.760 9.205 2.990 ;
        RECT  6.175 3.995 9.205 4.225 ;
        RECT  8.855 2.115 9.085 2.990 ;
        RECT  8.650 2.115 8.855 2.455 ;
        RECT  8.545 0.630 8.775 1.830 ;
        RECT  8.620 3.315 8.750 3.655 ;
        RECT  8.390 2.705 8.620 3.655 ;
        RECT  7.460 0.630 8.545 0.860 ;
        RECT  8.315 2.705 8.390 2.935 ;
        RECT  8.085 1.175 8.315 2.935 ;
        RECT  7.665 1.905 8.085 2.245 ;
        RECT  7.445 3.320 7.785 3.660 ;
        RECT  7.435 0.630 7.460 1.485 ;
        RECT  7.440 3.320 7.445 3.605 ;
        RECT  7.435 2.625 7.440 3.605 ;
        RECT  7.230 0.630 7.435 3.605 ;
        RECT  7.210 1.145 7.230 3.605 ;
        RECT  7.205 1.145 7.210 3.550 ;
        RECT  7.120 1.145 7.205 1.485 ;
        RECT  6.440 2.570 7.205 2.910 ;
        RECT  6.635 1.890 6.975 2.230 ;
        RECT  5.810 1.890 6.635 2.120 ;
        RECT  5.890 3.890 6.175 4.225 ;
        RECT  5.350 3.890 5.890 4.150 ;
        RECT  5.580 0.685 5.810 3.590 ;
        RECT  5.040 0.685 5.580 0.915 ;
        RECT  5.120 1.500 5.350 4.150 ;
        RECT  5.050 1.500 5.120 1.730 ;
        RECT  4.365 3.920 5.120 4.150 ;
        RECT  4.710 1.390 5.050 1.730 ;
        RECT  4.550 3.315 4.890 3.655 ;
        RECT  4.240 0.670 4.580 1.035 ;
        RECT  3.860 3.425 4.550 3.655 ;
        RECT  4.135 3.920 4.365 4.410 ;
        RECT  1.885 0.805 4.240 1.035 ;
        RECT  1.840 4.180 4.135 4.410 ;
        RECT  3.630 3.425 3.860 3.930 ;
        RECT  2.210 1.335 3.630 1.565 ;
        RECT  2.070 3.700 3.630 3.930 ;
        RECT  2.310 3.060 2.650 3.400 ;
        RECT  1.940 3.060 2.310 3.290 ;
        RECT  1.870 1.335 2.210 1.785 ;
        RECT  1.780 2.905 1.940 3.290 ;
        RECT  1.520 0.645 1.885 1.035 ;
        RECT  1.780 1.555 1.870 1.785 ;
        RECT  1.610 4.005 1.840 4.410 ;
        RECT  1.550 1.555 1.780 3.290 ;
        RECT  0.620 4.005 1.610 4.235 ;
        RECT  0.350 2.880 0.620 4.235 ;
        RECT  0.350 0.845 0.600 1.655 ;
        RECT  0.280 0.845 0.350 4.235 ;
        RECT  0.260 0.845 0.280 3.255 ;
        RECT  0.120 1.135 0.260 3.255 ;
    END
END SDFFX4

MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.870 1.820 3.160 2.100 ;
        RECT  2.520 1.730 2.870 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.055 2.720 4.165 3.060 ;
        RECT  3.825 2.405 4.055 3.060 ;
        RECT  3.820 2.405 3.825 2.660 ;
        RECT  2.500 2.405 3.820 2.635 ;
        RECT  2.050 2.380 2.500 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.395 1.355 15.625 3.330 ;
        RECT  15.320 1.355 15.395 1.845 ;
        RECT  15.340 3.100 15.395 3.330 ;
        RECT  15.000 3.100 15.340 3.440 ;
        RECT  15.220 1.355 15.320 1.695 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.860 0.700 14.200 1.080 ;
        RECT  13.505 0.850 13.860 1.080 ;
        RECT  13.720 2.870 13.800 3.210 ;
        RECT  13.505 2.380 13.720 3.210 ;
        RECT  13.460 0.850 13.505 3.210 ;
        RECT  13.340 0.850 13.460 2.660 ;
        RECT  13.275 0.850 13.340 2.610 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.965 1.405 4.465 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.150 1.235 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.320 -0.400 16.500 0.400 ;
        RECT  15.980 -0.400 16.320 0.575 ;
        RECT  15.000 -0.400 15.980 0.400 ;
        RECT  14.660 -0.400 15.000 0.575 ;
        RECT  13.400 -0.400 14.660 0.400 ;
        RECT  13.060 -0.400 13.400 0.575 ;
        RECT  11.440 -0.400 13.060 0.400 ;
        RECT  11.100 -0.400 11.440 1.270 ;
        RECT  8.825 -0.400 11.100 0.400 ;
        RECT  8.485 -0.400 8.825 1.445 ;
        RECT  6.660 -0.400 8.485 0.400 ;
        RECT  6.320 -0.400 6.660 1.270 ;
        RECT  3.140 -0.400 6.320 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.210 -0.400 2.800 0.400 ;
        RECT  1.210 1.440 1.240 1.780 ;
        RECT  0.870 -0.400 1.210 1.780 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.100 4.640 16.500 5.440 ;
        RECT  15.760 4.465 16.100 5.440 ;
        RECT  14.560 4.640 15.760 5.440 ;
        RECT  14.220 4.465 14.560 5.440 ;
        RECT  12.580 4.640 14.220 5.440 ;
        RECT  10.830 4.465 12.580 5.440 ;
        RECT  8.530 4.640 10.830 5.440 ;
        RECT  7.250 4.465 8.530 5.440 ;
        RECT  4.100 4.640 7.250 5.440 ;
        RECT  3.760 4.410 4.100 5.440 ;
        RECT  1.315 4.640 3.760 5.440 ;
        RECT  0.975 4.465 1.315 5.440 ;
        RECT  0.000 4.640 0.975 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.790 3.920 15.130 4.360 ;
        RECT  14.765 3.920 14.790 4.150 ;
        RECT  14.535 1.590 14.765 4.150 ;
        RECT  14.200 1.590 14.535 1.820 ;
        RECT  13.800 3.920 14.535 4.150 ;
        RECT  14.075 2.285 14.305 3.670 ;
        RECT  13.860 1.480 14.200 1.820 ;
        RECT  13.220 3.440 14.075 3.670 ;
        RECT  13.460 3.920 13.800 4.370 ;
        RECT  12.620 3.920 13.460 4.150 ;
        RECT  12.990 3.065 13.220 3.670 ;
        RECT  12.615 3.065 12.990 3.295 ;
        RECT  12.280 3.810 12.620 4.150 ;
        RECT  12.385 1.775 12.615 3.295 ;
        RECT  12.240 1.775 12.385 2.005 ;
        RECT  11.670 3.065 12.385 3.295 ;
        RECT  12.010 1.155 12.240 2.005 ;
        RECT  11.750 2.350 12.090 2.690 ;
        RECT  11.900 1.155 12.010 1.795 ;
        RECT  10.770 1.565 11.900 1.795 ;
        RECT  9.940 2.405 11.750 2.635 ;
        RECT  11.560 3.065 11.670 3.700 ;
        RECT  11.385 3.065 11.560 3.960 ;
        RECT  11.330 3.360 11.385 3.960 ;
        RECT  9.850 3.730 11.330 3.960 ;
        RECT  10.540 1.160 10.770 1.795 ;
        RECT  10.160 1.160 10.540 1.390 ;
        RECT  9.820 1.050 10.160 1.390 ;
        RECT  9.830 2.405 9.940 3.160 ;
        RECT  9.510 3.440 9.850 4.250 ;
        RECT  9.600 1.730 9.830 3.160 ;
        RECT  8.510 1.730 9.600 1.960 ;
        RECT  8.970 2.930 9.600 3.160 ;
        RECT  8.910 2.245 9.250 2.585 ;
        RECT  8.740 2.930 8.970 4.235 ;
        RECT  8.500 2.355 8.910 2.585 ;
        RECT  6.295 4.005 8.740 4.235 ;
        RECT  8.170 1.730 8.510 2.070 ;
        RECT  8.270 2.355 8.500 3.775 ;
        RECT  7.335 3.545 8.270 3.775 ;
        RECT  7.935 1.105 8.085 1.445 ;
        RECT  7.935 2.625 7.970 2.965 ;
        RECT  7.705 0.630 7.935 2.965 ;
        RECT  7.575 0.630 7.705 0.860 ;
        RECT  7.630 2.625 7.705 2.965 ;
        RECT  7.325 2.270 7.335 3.775 ;
        RECT  7.105 0.950 7.325 3.775 ;
        RECT  7.095 0.950 7.105 2.510 ;
        RECT  6.225 2.170 7.095 2.510 ;
        RECT  5.995 1.555 6.820 1.785 ;
        RECT  6.290 3.890 6.295 4.235 ;
        RECT  5.950 3.890 6.290 4.280 ;
        RECT  5.765 1.545 5.995 3.600 ;
        RECT  5.535 3.890 5.950 4.150 ;
        RECT  5.610 1.545 5.765 1.785 ;
        RECT  5.380 0.920 5.610 1.785 ;
        RECT  5.305 2.765 5.535 4.150 ;
        RECT  5.300 0.920 5.380 1.150 ;
        RECT  5.070 2.765 5.305 2.995 ;
        RECT  3.530 3.920 5.305 4.150 ;
        RECT  4.960 0.810 5.300 1.150 ;
        RECT  4.735 3.260 5.075 3.600 ;
        RECT  4.840 1.380 5.070 2.995 ;
        RECT  4.730 1.380 4.840 1.720 ;
        RECT  3.070 3.370 4.735 3.600 ;
        RECT  4.160 0.750 4.500 1.090 ;
        RECT  2.555 0.810 4.160 1.040 ;
        RECT  3.210 1.270 3.550 1.575 ;
        RECT  3.300 3.920 3.530 4.410 ;
        RECT  1.980 4.180 3.300 4.410 ;
        RECT  2.120 1.270 3.210 1.500 ;
        RECT  2.840 3.370 3.070 3.930 ;
        RECT  2.295 3.700 2.840 3.930 ;
        RECT  2.270 3.040 2.610 3.380 ;
        RECT  2.325 0.645 2.555 1.040 ;
        RECT  1.440 0.645 2.325 0.875 ;
        RECT  2.080 3.040 2.270 3.270 ;
        RECT  1.835 1.270 2.120 1.780 ;
        RECT  1.820 2.940 2.080 3.270 ;
        RECT  1.750 3.605 1.980 4.410 ;
        RECT  1.820 1.440 1.835 1.780 ;
        RECT  1.780 1.440 1.820 3.270 ;
        RECT  1.590 1.550 1.780 3.270 ;
        RECT  0.570 3.605 1.750 3.835 ;
        RECT  0.340 1.340 0.570 3.835 ;
        RECT  0.180 1.340 0.340 1.680 ;
        RECT  0.180 3.025 0.340 3.365 ;
    END
END SDFFX2

MACRO SDFFX1
    CLASS CORE ;
    FOREIGN SDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.845 3.290 2.380 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 2.630 3.615 3.030 ;
        RECT  2.500 2.630 3.275 2.860 ;
        RECT  2.210 2.380 2.500 2.860 ;
        RECT  2.120 2.380 2.210 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.340 1.190 13.680 3.880 ;
        RECT  13.240 3.540 13.340 3.880 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 0.865 12.985 3.420 ;
        RECT  12.285 0.865 12.755 1.095 ;
        RECT  11.870 3.190 12.755 3.420 ;
        RECT  11.940 0.695 12.285 1.095 ;
        RECT  11.530 3.190 11.870 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 1.845 4.405 2.075 ;
        RECT  4.015 1.405 4.270 2.075 ;
        RECT  3.930 1.405 4.015 1.745 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.205 1.180 2.660 ;
        RECT  0.645 2.150 0.875 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 -0.400 13.860 0.400 ;
        RECT  12.680 -0.400 13.020 0.575 ;
        RECT  11.520 -0.400 12.680 0.400 ;
        RECT  11.180 -0.400 11.520 0.575 ;
        RECT  9.080 -0.400 11.180 0.400 ;
        RECT  8.740 -0.400 9.080 1.460 ;
        RECT  6.710 -0.400 8.740 0.400 ;
        RECT  6.370 -0.400 6.710 1.150 ;
        RECT  3.190 -0.400 6.370 0.400 ;
        RECT  2.850 -0.400 3.190 0.575 ;
        RECT  1.260 -0.400 2.850 0.400 ;
        RECT  1.260 1.345 1.510 1.685 ;
        RECT  1.030 -0.400 1.260 1.685 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.630 4.640 13.860 5.440 ;
        RECT  12.290 4.410 12.630 5.440 ;
        RECT  11.110 4.640 12.290 5.440 ;
        RECT  10.770 4.465 11.110 5.440 ;
        RECT  8.435 4.640 10.770 5.440 ;
        RECT  8.095 4.465 8.435 5.440 ;
        RECT  6.925 4.640 8.095 5.440 ;
        RECT  6.585 4.465 6.925 5.440 ;
        RECT  3.885 4.640 6.585 5.440 ;
        RECT  3.545 4.410 3.885 5.440 ;
        RECT  1.100 4.640 3.545 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.450 1.470 12.510 2.350 ;
        RECT  12.280 1.470 12.450 2.900 ;
        RECT  11.980 1.470 12.280 1.810 ;
        RECT  12.220 2.120 12.280 2.900 ;
        RECT  11.040 2.670 12.220 2.900 ;
        RECT  11.555 2.045 11.895 2.385 ;
        RECT  11.760 4.065 11.870 4.405 ;
        RECT  11.530 3.970 11.760 4.405 ;
        RECT  11.520 2.045 11.555 2.275 ;
        RECT  11.040 3.970 11.530 4.200 ;
        RECT  11.290 1.550 11.520 2.275 ;
        RECT  10.360 1.550 11.290 1.780 ;
        RECT  10.810 2.180 11.040 4.200 ;
        RECT  10.650 2.180 10.810 2.520 ;
        RECT  10.400 0.820 10.740 1.160 ;
        RECT  9.580 0.930 10.400 1.160 ;
        RECT  10.190 1.440 10.360 1.780 ;
        RECT  9.960 1.440 10.190 4.010 ;
        RECT  9.850 3.780 9.960 4.010 ;
        RECT  9.510 3.780 9.850 4.120 ;
        RECT  9.580 2.820 9.730 3.160 ;
        RECT  9.350 0.930 9.580 3.515 ;
        RECT  8.200 1.755 9.350 1.985 ;
        RECT  8.910 3.285 9.350 3.515 ;
        RECT  8.720 2.370 9.060 2.710 ;
        RECT  8.680 3.285 8.910 4.235 ;
        RECT  8.440 2.480 8.720 2.710 ;
        RECT  5.845 4.005 8.680 4.235 ;
        RECT  8.210 2.480 8.440 3.775 ;
        RECT  8.100 1.170 8.250 1.510 ;
        RECT  7.075 3.545 8.210 3.775 ;
        RECT  7.955 0.630 8.100 1.510 ;
        RECT  7.755 0.630 7.955 3.075 ;
        RECT  7.725 0.630 7.755 3.130 ;
        RECT  7.415 2.790 7.725 3.130 ;
        RECT  7.225 0.810 7.455 2.470 ;
        RECT  7.075 2.130 7.225 2.470 ;
        RECT  6.845 2.130 7.075 3.775 ;
        RECT  6.655 1.460 6.995 1.800 ;
        RECT  6.090 2.130 6.845 2.470 ;
        RECT  5.550 1.570 6.655 1.800 ;
        RECT  5.505 3.950 5.845 4.290 ;
        RECT  5.320 0.745 5.550 3.680 ;
        RECT  5.085 3.950 5.505 4.180 ;
        RECT  5.065 0.745 5.320 1.090 ;
        RECT  4.855 1.340 5.085 4.180 ;
        RECT  5.010 0.750 5.065 1.090 ;
        RECT  4.730 1.340 4.855 1.680 ;
        RECT  3.315 3.950 4.855 4.180 ;
        RECT  2.855 3.320 4.625 3.660 ;
        RECT  4.210 0.750 4.550 1.090 ;
        RECT  2.605 0.810 4.210 1.040 ;
        RECT  2.310 1.345 3.595 1.575 ;
        RECT  3.085 3.950 3.315 4.410 ;
        RECT  1.565 4.180 3.085 4.410 ;
        RECT  2.625 3.320 2.855 3.930 ;
        RECT  1.800 3.700 2.625 3.930 ;
        RECT  2.375 0.645 2.605 1.040 ;
        RECT  1.890 3.095 2.395 3.325 ;
        RECT  1.490 0.645 2.375 0.875 ;
        RECT  2.025 1.345 2.310 1.770 ;
        RECT  1.970 1.430 2.025 1.770 ;
        RECT  1.890 1.540 1.970 2.145 ;
        RECT  1.740 1.540 1.890 3.325 ;
        RECT  1.660 1.915 1.740 3.325 ;
        RECT  1.520 2.885 1.660 3.325 ;
        RECT  1.335 3.605 1.565 4.410 ;
        RECT  0.570 3.605 1.335 3.835 ;
        RECT  0.410 1.430 0.750 1.770 ;
        RECT  0.380 3.020 0.570 3.835 ;
        RECT  0.380 1.540 0.410 1.770 ;
        RECT  0.150 1.540 0.380 3.835 ;
    END
END SDFFX1

MACRO RSLATNXL
    CLASS CORE ;
    FOREIGN RSLATNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.290 1.845 2.835 2.450 ;
        RECT  2.195 1.845 2.290 2.075 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.415 2.270 3.855 2.820 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.100 6.335 3.755 ;
        RECT  5.495 2.965 6.105 3.195 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 3.545 0.520 3.885 ;
        RECT  0.410 1.100 0.465 1.450 ;
        RECT  0.410 3.525 0.465 3.885 ;
        RECT  0.180 1.100 0.410 3.885 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 -0.400 6.600 0.400 ;
        RECT  5.380 -0.400 5.720 0.575 ;
        RECT  4.215 -0.400 5.380 0.400 ;
        RECT  3.875 -0.400 4.215 0.575 ;
        RECT  2.800 -0.400 3.875 0.400 ;
        RECT  2.460 -0.400 2.800 0.575 ;
        RECT  1.080 -0.400 2.460 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.560 4.640 6.600 5.440 ;
        RECT  5.220 4.465 5.560 5.440 ;
        RECT  2.610 4.640 5.220 5.440 ;
        RECT  2.270 4.465 2.610 5.440 ;
        RECT  1.240 4.640 2.270 5.440 ;
        RECT  0.900 3.765 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.625 0.870 5.855 2.655 ;
        RECT  4.965 0.870 5.625 1.100 ;
        RECT  4.920 2.255 5.625 2.485 ;
        RECT  4.790 1.640 5.300 1.870 ;
        RECT  4.735 0.750 4.965 1.100 ;
        RECT  4.690 2.255 4.920 3.840 ;
        RECT  4.560 1.335 4.790 1.870 ;
        RECT  4.140 3.610 4.690 3.840 ;
        RECT  4.490 1.335 4.560 1.565 ;
        RECT  4.260 0.805 4.490 1.565 ;
        RECT  4.090 1.805 4.320 3.375 ;
        RECT  1.905 0.805 4.260 1.035 ;
        RECT  3.910 3.610 4.140 4.410 ;
        RECT  4.030 1.805 4.090 2.035 ;
        RECT  3.680 3.145 4.090 3.375 ;
        RECT  3.800 1.330 4.030 2.035 ;
        RECT  3.080 4.180 3.910 4.410 ;
        RECT  3.450 3.145 3.680 3.845 ;
        RECT  1.740 2.760 3.170 2.990 ;
        RECT  2.850 4.000 3.080 4.410 ;
        RECT  1.740 4.000 2.850 4.230 ;
        RECT  1.740 1.265 2.680 1.495 ;
        RECT  1.540 0.665 1.905 1.035 ;
        RECT  1.510 1.265 1.740 2.990 ;
        RECT  0.930 0.805 1.540 1.035 ;
        RECT  1.325 1.580 1.510 1.945 ;
        RECT  0.930 2.900 1.280 3.130 ;
        RECT  0.700 0.805 0.930 3.130 ;
        RECT  0.645 2.100 0.700 2.475 ;
    END
END RSLATNXL

MACRO RSLATNX4
    CLASS CORE ;
    FOREIGN RSLATNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATNXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 1.845 2.155 2.490 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 1.685 9.760 2.280 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.770 0.920 10.880 1.730 ;
        RECT  10.755 0.920 10.770 2.635 ;
        RECT  10.540 0.920 10.755 3.090 ;
        RECT  10.420 1.820 10.540 3.090 ;
        RECT  10.040 1.820 10.420 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 2.635 1.240 3.035 ;
        RECT  0.875 1.260 1.180 3.035 ;
        RECT  0.800 1.260 0.875 2.660 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.600 -0.400 11.880 0.400 ;
        RECT  11.260 -0.400 11.600 1.425 ;
        RECT  10.160 -0.400 11.260 0.400 ;
        RECT  9.820 -0.400 10.160 1.295 ;
        RECT  8.810 -0.400 9.820 0.400 ;
        RECT  8.470 -0.400 8.810 0.575 ;
        RECT  7.450 -0.400 8.470 0.400 ;
        RECT  7.110 -0.400 7.450 0.950 ;
        RECT  6.090 -0.400 7.110 0.400 ;
        RECT  5.750 -0.400 6.090 0.950 ;
        RECT  4.725 -0.400 5.750 0.400 ;
        RECT  4.385 -0.400 4.725 0.950 ;
        RECT  3.360 -0.400 4.385 0.400 ;
        RECT  3.020 -0.400 3.360 0.575 ;
        RECT  1.800 -0.400 3.020 0.400 ;
        RECT  1.460 -0.400 1.800 0.965 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.965 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.530 4.640 11.880 5.440 ;
        RECT  11.190 4.090 11.530 5.440 ;
        RECT  10.090 4.640 11.190 5.440 ;
        RECT  9.750 4.090 10.090 5.440 ;
        RECT  8.580 4.640 9.750 5.440 ;
        RECT  8.240 4.090 8.580 5.440 ;
        RECT  6.020 4.640 8.240 5.440 ;
        RECT  5.680 3.620 6.020 5.440 ;
        RECT  3.260 4.640 5.680 5.440 ;
        RECT  2.920 3.795 3.260 5.440 ;
        RECT  1.960 4.640 2.920 5.440 ;
        RECT  1.620 3.735 1.960 5.440 ;
        RECT  0.520 4.640 1.620 5.440 ;
        RECT  0.180 4.090 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.005 2.210 11.235 3.685 ;
        RECT  8.615 3.455 11.005 3.685 ;
        RECT  9.075 1.090 9.435 1.320 ;
        RECT  9.075 2.805 9.325 3.035 ;
        RECT  8.845 1.090 9.075 3.035 ;
        RECT  8.385 1.210 8.615 3.685 ;
        RECT  8.130 1.210 8.385 1.440 ;
        RECT  7.300 3.455 8.385 3.685 ;
        RECT  7.925 2.110 8.155 2.500 ;
        RECT  7.790 1.155 8.130 1.495 ;
        RECT  5.740 2.270 7.925 2.500 ;
        RECT  6.770 1.210 7.790 1.440 ;
        RECT  6.960 2.835 7.300 4.115 ;
        RECT  6.430 1.155 6.770 1.495 ;
        RECT  6.040 1.210 6.430 1.440 ;
        RECT  5.810 1.210 6.040 2.040 ;
        RECT  3.775 1.810 5.810 2.040 ;
        RECT  5.510 2.270 5.740 3.065 ;
        RECT  4.740 2.835 5.510 3.065 ;
        RECT  5.065 1.155 5.405 1.495 ;
        RECT  4.045 1.210 5.065 1.440 ;
        RECT  4.400 2.835 4.740 4.115 ;
        RECT  3.315 3.235 4.400 3.500 ;
        RECT  3.705 1.155 4.045 1.495 ;
        RECT  3.545 1.810 3.775 2.555 ;
        RECT  3.315 1.210 3.705 1.440 ;
        RECT  3.085 1.210 3.315 3.500 ;
        RECT  0.570 3.270 3.085 3.500 ;
        RECT  2.625 1.270 2.855 3.035 ;
        RECT  2.220 1.270 2.625 1.500 ;
        RECT  2.380 2.805 2.625 3.035 ;
        RECT  0.340 2.210 0.570 3.500 ;
    END
END RSLATNX4

MACRO RSLATNX2
    CLASS CORE ;
    FOREIGN RSLATNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATNXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 2.330 3.745 2.635 ;
        RECT  3.145 2.330 3.515 2.560 ;
        RECT  2.915 2.200 3.145 2.560 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.710 1.820 4.480 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.000 2.955 7.045 3.205 ;
        RECT  6.935 1.030 7.000 3.205 ;
        RECT  6.770 1.030 6.935 3.690 ;
        RECT  6.595 1.030 6.770 1.370 ;
        RECT  6.595 2.750 6.770 3.690 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.395 0.920 0.520 1.260 ;
        RECT  0.465 2.750 0.520 3.690 ;
        RECT  0.395 2.750 0.465 3.755 ;
        RECT  0.165 0.920 0.395 3.755 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.170 -0.400 7.260 0.400 ;
        RECT  5.830 -0.400 6.170 0.575 ;
        RECT  4.550 -0.400 5.830 0.400 ;
        RECT  4.210 -0.400 4.550 0.575 ;
        RECT  2.680 -0.400 4.210 0.400 ;
        RECT  2.340 -0.400 2.680 1.275 ;
        RECT  1.240 -0.400 2.340 0.400 ;
        RECT  0.900 -0.400 1.240 1.300 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.215 4.640 7.260 5.440 ;
        RECT  5.875 4.090 6.215 5.440 ;
        RECT  3.820 4.640 5.875 5.440 ;
        RECT  3.480 4.410 3.820 5.440 ;
        RECT  1.240 4.640 3.480 5.440 ;
        RECT  0.900 4.090 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.305 1.725 6.535 2.340 ;
        RECT  5.430 1.725 6.305 1.955 ;
        RECT  5.640 2.215 5.865 3.850 ;
        RECT  5.635 2.215 5.640 4.405 ;
        RECT  5.410 3.620 5.635 4.405 ;
        RECT  5.405 0.900 5.430 1.955 ;
        RECT  4.365 4.175 5.410 4.405 ;
        RECT  5.175 0.900 5.405 3.345 ;
        RECT  5.070 0.900 5.175 1.130 ;
        RECT  4.945 3.115 5.175 3.345 ;
        RECT  4.715 3.115 4.945 3.945 ;
        RECT  4.710 1.360 4.940 2.560 ;
        RECT  4.595 3.305 4.715 3.945 ;
        RECT  3.900 1.360 4.710 1.590 ;
        RECT  4.330 2.330 4.710 2.560 ;
        RECT  2.165 3.305 4.595 3.535 ;
        RECT  4.135 3.775 4.365 4.405 ;
        RECT  4.100 2.330 4.330 3.075 ;
        RECT  1.700 3.775 4.135 4.005 ;
        RECT  3.670 0.670 3.900 1.590 ;
        RECT  3.315 0.670 3.670 0.900 ;
        RECT  3.100 1.415 3.440 1.755 ;
        RECT  2.635 1.525 3.100 1.755 ;
        RECT  2.635 2.790 3.060 3.020 ;
        RECT  2.405 1.525 2.635 3.020 ;
        RECT  1.940 2.255 2.405 2.485 ;
        RECT  1.935 2.855 2.165 3.535 ;
        RECT  1.620 1.415 1.960 1.865 ;
        RECT  1.525 2.855 1.935 3.085 ;
        RECT  1.470 3.375 1.700 4.005 ;
        RECT  0.855 1.635 1.620 1.865 ;
        RECT  1.295 2.200 1.525 3.085 ;
        RECT  0.980 3.375 1.470 3.605 ;
        RECT  0.855 2.285 0.980 3.605 ;
        RECT  0.750 1.635 0.855 3.605 ;
        RECT  0.625 1.635 0.750 2.515 ;
    END
END RSLATNX2

MACRO RSLATNX1
    CLASS CORE ;
    FOREIGN RSLATNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATNXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.380 3.205 2.865 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.380 4.160 2.865 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.840 1.240 7.070 3.500 ;
        RECT  6.680 1.240 6.840 1.580 ;
        RECT  6.815 1.845 6.840 2.075 ;
        RECT  6.680 3.160 6.840 3.500 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.235 1.240 0.465 3.755 ;
        RECT  0.175 3.195 0.235 3.755 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.460 -0.400 7.260 0.400 ;
        RECT  6.120 -0.400 6.460 0.575 ;
        RECT  4.860 -0.400 6.120 0.400 ;
        RECT  4.520 -0.400 4.860 0.575 ;
        RECT  2.735 -0.400 4.520 0.400 ;
        RECT  2.395 -0.400 2.735 0.575 ;
        RECT  1.095 -0.400 2.395 0.400 ;
        RECT  0.755 -0.400 1.095 0.575 ;
        RECT  0.000 -0.400 0.755 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.460 4.640 7.260 5.440 ;
        RECT  6.120 4.465 6.460 5.440 ;
        RECT  3.595 4.640 6.120 5.440 ;
        RECT  3.255 4.465 3.595 5.440 ;
        RECT  1.240 4.640 3.255 5.440 ;
        RECT  0.900 3.765 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.350 2.685 6.610 2.915 ;
        RECT  6.120 0.870 6.350 2.915 ;
        RECT  5.320 0.870 6.120 1.100 ;
        RECT  5.795 2.685 6.120 2.915 ;
        RECT  5.655 1.335 5.885 2.400 ;
        RECT  5.565 2.685 5.795 4.050 ;
        RECT  4.420 1.335 5.655 1.565 ;
        RECT  2.890 3.820 5.565 4.050 ;
        RECT  5.095 1.855 5.325 3.350 ;
        RECT  3.960 1.855 5.095 2.085 ;
        RECT  4.260 3.120 5.095 3.350 ;
        RECT  4.190 0.805 4.420 1.565 ;
        RECT  1.890 0.805 4.190 1.035 ;
        RECT  3.730 1.350 3.960 2.085 ;
        RECT  2.365 3.115 3.800 3.345 ;
        RECT  2.660 3.820 2.890 4.375 ;
        RECT  2.355 4.145 2.660 4.375 ;
        RECT  2.365 1.405 2.615 1.635 ;
        RECT  2.135 1.405 2.365 3.345 ;
        RECT  1.560 1.405 2.135 1.635 ;
        RECT  1.515 0.700 1.890 1.035 ;
        RECT  1.500 2.825 1.730 3.400 ;
        RECT  1.330 1.405 1.560 1.765 ;
        RECT  0.945 0.805 1.515 1.035 ;
        RECT  0.945 2.825 1.500 3.055 ;
        RECT  0.715 0.805 0.945 3.055 ;
    END
END RSLATNX1

MACRO RSLATXL
    CLASS CORE ;
    FOREIGN RSLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.815 3.160 2.095 ;
        RECT  2.780 1.815 2.970 2.305 ;
        RECT  2.550 1.840 2.780 2.305 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.230 2.330 3.820 2.680 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.060 0.520 1.400 ;
        RECT  0.360 2.920 0.520 3.260 ;
        RECT  0.130 1.060 0.360 3.260 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.935 1.095 6.275 1.435 ;
        RECT  5.910 1.205 5.935 1.435 ;
        RECT  5.850 1.205 5.910 3.750 ;
        RECT  5.680 1.205 5.850 3.860 ;
        RECT  5.510 3.520 5.680 3.860 ;
        RECT  5.495 3.520 5.510 3.805 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.710 -0.400 6.600 0.400 ;
        RECT  5.370 -0.400 5.710 0.575 ;
        RECT  3.150 -0.400 5.370 0.400 ;
        RECT  2.810 -0.400 3.150 0.575 ;
        RECT  1.080 -0.400 2.810 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.090 4.640 6.600 5.440 ;
        RECT  4.750 4.465 5.090 5.440 ;
        RECT  1.750 4.640 4.750 5.440 ;
        RECT  0.940 4.465 1.750 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.745 2.330 5.445 2.670 ;
        RECT  4.515 0.835 4.745 3.860 ;
        RECT  4.350 0.835 4.515 1.065 ;
        RECT  4.190 3.520 4.515 3.860 ;
        RECT  4.010 0.725 4.350 1.065 ;
        RECT  4.050 1.540 4.280 3.290 ;
        RECT  4.095 3.630 4.190 3.860 ;
        RECT  3.865 3.630 4.095 4.410 ;
        RECT  3.850 1.540 4.050 1.770 ;
        RECT  3.635 3.060 4.050 3.290 ;
        RECT  2.220 4.180 3.865 4.410 ;
        RECT  3.510 1.430 3.850 1.770 ;
        RECT  3.380 0.630 3.720 1.035 ;
        RECT  3.405 3.060 3.635 3.945 ;
        RECT  2.870 3.715 3.405 3.945 ;
        RECT  2.525 0.805 3.380 1.035 ;
        RECT  2.830 2.920 3.170 3.260 ;
        RECT  2.315 2.920 2.830 3.150 ;
        RECT  2.295 0.665 2.525 1.035 ;
        RECT  2.315 1.365 2.450 1.595 ;
        RECT  2.085 1.365 2.315 3.150 ;
        RECT  1.665 0.665 2.295 0.895 ;
        RECT  1.990 3.870 2.220 4.410 ;
        RECT  1.750 2.340 2.085 2.680 ;
        RECT  1.610 3.870 1.990 4.100 ;
        RECT  1.510 2.920 1.850 3.260 ;
        RECT  1.435 0.665 1.665 1.205 ;
        RECT  1.270 3.760 1.610 4.100 ;
        RECT  1.025 2.975 1.510 3.205 ;
        RECT  1.025 0.975 1.435 1.205 ;
        RECT  0.795 0.975 1.025 3.205 ;
        RECT  0.590 1.790 0.795 2.130 ;
    END
END RSLATXL

MACRO RSLATX4
    CLASS CORE ;
    FOREIGN RSLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.195 1.845 9.760 2.240 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.725 2.205 2.500 2.660 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.420 1.325 10.645 1.665 ;
        RECT  10.420 2.875 10.540 3.215 ;
        RECT  10.190 1.325 10.420 3.220 ;
        RECT  10.040 1.820 10.190 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 1.820 1.180 3.220 ;
        RECT  0.820 1.325 1.160 3.220 ;
        RECT  0.800 1.820 0.820 3.220 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.285 -0.400 11.880 0.400 ;
        RECT  10.945 -0.400 11.285 0.955 ;
        RECT  10.005 -0.400 10.945 0.400 ;
        RECT  9.665 -0.400 10.005 0.955 ;
        RECT  8.730 -0.400 9.665 0.400 ;
        RECT  8.390 -0.400 8.730 0.575 ;
        RECT  6.130 -0.400 8.390 0.400 ;
        RECT  5.790 -0.400 6.130 0.955 ;
        RECT  3.460 -0.400 5.790 0.400 ;
        RECT  3.120 -0.400 3.460 1.135 ;
        RECT  1.800 -0.400 3.120 0.400 ;
        RECT  1.460 -0.400 1.800 0.965 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.965 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.180 4.640 11.880 5.440 ;
        RECT  10.840 4.145 11.180 5.440 ;
        RECT  9.900 4.640 10.840 5.440 ;
        RECT  9.560 4.145 9.900 5.440 ;
        RECT  8.520 4.640 9.560 5.440 ;
        RECT  8.180 4.465 8.520 5.440 ;
        RECT  7.200 4.640 8.180 5.440 ;
        RECT  6.860 3.765 7.200 5.440 ;
        RECT  5.920 4.640 6.860 5.440 ;
        RECT  5.580 3.765 5.920 5.440 ;
        RECT  4.635 4.640 5.580 5.440 ;
        RECT  4.295 3.765 4.635 5.440 ;
        RECT  3.270 4.640 4.295 5.440 ;
        RECT  2.930 4.465 3.270 5.440 ;
        RECT  1.800 4.640 2.930 5.440 ;
        RECT  1.460 4.145 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 4.145 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.770 2.210 11.000 3.895 ;
        RECT  8.110 3.665 10.770 3.895 ;
        RECT  8.895 1.360 9.235 1.590 ;
        RECT  8.895 3.155 9.115 3.385 ;
        RECT  8.665 1.360 8.895 3.385 ;
        RECT  7.820 1.915 8.325 2.145 ;
        RECT  7.880 2.975 8.110 3.895 ;
        RECT  7.355 2.975 7.880 3.205 ;
        RECT  7.590 0.855 7.820 2.145 ;
        RECT  6.690 0.855 7.590 1.085 ;
        RECT  7.125 1.315 7.355 3.205 ;
        RECT  5.750 2.975 7.125 3.205 ;
        RECT  6.460 0.855 6.690 1.600 ;
        RECT  6.265 1.370 6.460 1.600 ;
        RECT  6.035 1.370 6.265 2.725 ;
        RECT  4.795 1.370 6.035 1.600 ;
        RECT  5.520 2.445 5.750 3.205 ;
        RECT  3.885 2.445 5.520 2.675 ;
        RECT  3.425 2.975 5.280 3.205 ;
        RECT  4.510 1.365 4.795 1.600 ;
        RECT  3.425 1.365 4.510 1.595 ;
        RECT  3.655 1.860 3.885 2.675 ;
        RECT  3.195 1.365 3.425 3.910 ;
        RECT  0.495 3.680 3.195 3.910 ;
        RECT  2.730 1.420 2.960 3.445 ;
        RECT  2.225 1.420 2.730 1.650 ;
        RECT  2.225 3.215 2.730 3.445 ;
        RECT  0.265 2.210 0.495 3.910 ;
    END
END RSLATX4

MACRO RSLATX2
    CLASS CORE ;
    FOREIGN RSLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.585 2.035 6.385 2.635 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.795 1.560 3.255 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.545 0.940 7.600 1.845 ;
        RECT  7.315 0.940 7.545 3.125 ;
        RECT  7.260 0.940 7.315 1.750 ;
        RECT  7.045 2.895 7.315 3.125 ;
        RECT  7.010 2.895 7.045 3.195 ;
        RECT  6.670 2.895 7.010 4.175 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 0.790 0.520 1.730 ;
        RECT  0.360 2.750 0.520 4.030 ;
        RECT  0.180 0.790 0.360 4.030 ;
        RECT  0.130 0.790 0.180 2.985 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.835 -0.400 7.920 0.400 ;
        RECT  6.495 -0.400 6.835 0.575 ;
        RECT  4.255 -0.400 6.495 0.400 ;
        RECT  3.915 -0.400 4.255 0.575 ;
        RECT  2.040 -0.400 3.915 0.400 ;
        RECT  1.230 -0.400 2.040 0.575 ;
        RECT  0.000 -0.400 1.230 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.215 4.640 7.920 5.440 ;
        RECT  5.875 4.090 6.215 5.440 ;
        RECT  5.165 4.640 5.875 5.440 ;
        RECT  4.825 3.635 5.165 5.440 ;
        RECT  3.670 4.640 4.825 5.440 ;
        RECT  3.330 4.465 3.670 5.440 ;
        RECT  2.550 4.640 3.330 5.440 ;
        RECT  2.210 4.465 2.550 5.440 ;
        RECT  1.280 4.640 2.210 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.010 2.220 7.065 2.560 ;
        RECT  6.780 0.805 7.010 2.560 ;
        RECT  5.575 0.805 6.780 1.035 ;
        RECT  6.725 2.220 6.780 2.560 ;
        RECT  5.775 1.450 6.115 1.790 ;
        RECT  5.155 1.505 5.775 1.735 ;
        RECT  5.350 2.890 5.690 3.230 ;
        RECT  5.235 0.750 5.575 1.090 ;
        RECT  5.155 2.890 5.350 3.120 ;
        RECT  4.595 0.805 5.235 1.035 ;
        RECT  5.155 2.215 5.210 2.555 ;
        RECT  4.925 1.505 5.155 3.120 ;
        RECT  4.870 2.215 4.925 2.555 ;
        RECT  4.365 0.805 4.595 3.875 ;
        RECT  4.090 3.510 4.365 3.875 ;
        RECT  3.905 1.240 4.135 3.175 ;
        RECT  2.485 3.645 4.090 3.875 ;
        RECT  3.710 1.240 3.905 1.470 ;
        RECT  3.110 2.945 3.905 3.175 ;
        RECT  3.605 1.130 3.710 1.470 ;
        RECT  3.370 0.920 3.605 1.470 ;
        RECT  3.130 1.860 3.470 2.200 ;
        RECT  0.980 0.920 3.370 1.150 ;
        RECT  3.060 1.860 3.130 2.090 ;
        RECT  2.770 2.945 3.110 3.285 ;
        RECT  2.830 1.445 3.060 2.090 ;
        RECT  2.020 1.445 2.830 1.675 ;
        RECT  2.485 2.200 2.595 2.540 ;
        RECT  2.255 2.200 2.485 3.875 ;
        RECT  1.890 1.445 2.020 3.920 ;
        RECT  1.790 1.390 1.890 3.920 ;
        RECT  1.550 1.390 1.790 1.730 ;
        RECT  1.510 3.580 1.790 3.920 ;
        RECT  0.750 0.920 0.980 2.365 ;
        RECT  0.600 2.025 0.750 2.365 ;
    END
END RSLATX2

MACRO RSLATX1
    CLASS CORE ;
    FOREIGN RSLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.880 1.820 3.160 2.100 ;
        RECT  2.650 1.820 2.880 2.565 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.115 2.330 3.820 2.720 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.240 0.520 1.580 ;
        RECT  0.405 2.955 0.520 3.295 ;
        RECT  0.175 1.240 0.405 3.295 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.155 1.190 6.310 1.530 ;
        RECT  5.970 1.190 6.155 1.540 ;
        RECT  5.855 1.300 5.970 1.540 ;
        RECT  5.855 3.545 5.915 3.885 ;
        RECT  5.625 1.300 5.855 3.885 ;
        RECT  5.575 3.525 5.625 3.885 ;
        RECT  5.495 3.525 5.575 3.830 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.745 -0.400 6.600 0.400 ;
        RECT  5.405 -0.400 5.745 0.575 ;
        RECT  3.160 -0.400 5.405 0.400 ;
        RECT  2.820 -0.400 3.160 0.575 ;
        RECT  1.085 -0.400 2.820 0.400 ;
        RECT  0.745 -0.400 1.085 0.575 ;
        RECT  0.000 -0.400 0.745 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 4.640 6.600 5.440 ;
        RECT  4.760 4.465 5.100 5.440 ;
        RECT  1.755 4.640 4.760 5.440 ;
        RECT  0.945 4.465 1.755 5.440 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.165 1.000 5.395 3.065 ;
        RECT  4.415 1.000 5.165 1.230 ;
        RECT  4.750 2.835 5.165 3.065 ;
        RECT  4.520 2.835 4.750 3.860 ;
        RECT  4.335 3.520 4.520 3.860 ;
        RECT  4.075 0.945 4.415 1.285 ;
        RECT  4.105 3.520 4.335 4.405 ;
        RECT  4.055 1.755 4.285 3.290 ;
        RECT  2.645 4.175 4.105 4.405 ;
        RECT  3.885 1.755 4.055 1.985 ;
        RECT  3.660 3.060 4.055 3.290 ;
        RECT  3.545 1.645 3.885 1.985 ;
        RECT  3.440 0.810 3.780 1.150 ;
        RECT  3.430 3.060 3.660 3.940 ;
        RECT  2.415 0.865 3.440 1.095 ;
        RECT  2.875 3.710 3.430 3.940 ;
        RECT  2.835 2.955 3.175 3.295 ;
        RECT  2.400 2.955 2.835 3.185 ;
        RECT  2.415 3.810 2.645 4.405 ;
        RECT  2.075 0.750 2.415 1.095 ;
        RECT  1.615 3.810 2.415 4.040 ;
        RECT  2.170 1.450 2.400 3.185 ;
        RECT  1.835 2.110 2.170 2.450 ;
        RECT  1.100 0.865 2.075 1.095 ;
        RECT  1.515 3.075 1.855 3.415 ;
        RECT  1.275 3.755 1.615 4.095 ;
        RECT  1.100 3.130 1.515 3.360 ;
        RECT  0.870 0.865 1.100 3.360 ;
        RECT  0.640 1.905 0.870 2.270 ;
    END
END RSLATX1

MACRO OR4XL
    CLASS CORE ;
    FOREIGN OR4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.060 3.820 3.870 ;
        RECT  3.420 1.060 3.590 1.400 ;
        RECT  3.440 3.195 3.590 3.870 ;
        RECT  3.240 3.365 3.440 3.870 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.715 2.330 3.190 2.795 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 2.330 1.980 3.220 ;
        RECT  1.460 2.910 1.750 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.170 1.280 2.665 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.755 0.560 3.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.000 -0.400 3.960 0.400 ;
        RECT  2.660 -0.400 3.000 0.575 ;
        RECT  1.120 -0.400 2.660 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.245 4.640 3.960 5.440 ;
        RECT  2.435 4.465 3.245 5.440 ;
        RECT  0.000 4.640 2.435 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.480 1.655 3.295 2.005 ;
        RECT  2.250 1.180 2.480 3.915 ;
        RECT  2.060 1.180 2.250 1.520 ;
        RECT  0.540 3.685 2.250 3.915 ;
        RECT  0.800 1.180 2.060 1.410 ;
        RECT  0.570 1.180 0.800 1.780 ;
        RECT  0.460 1.440 0.570 1.780 ;
        RECT  0.200 3.630 0.540 3.970 ;
    END
END OR4XL

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR4XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 1.445 6.080 3.330 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 1.740 4.955 3.730 ;
        RECT  4.615 1.740 4.725 1.970 ;
        RECT  1.540 3.500 4.725 3.730 ;
        RECT  4.275 1.630 4.615 1.970 ;
        RECT  0.800 3.500 1.540 3.890 ;
        RECT  0.700 3.500 0.800 3.755 ;
        RECT  0.470 2.605 0.700 3.755 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 2.300 4.435 2.640 ;
        RECT  4.150 2.300 4.380 3.260 ;
        RECT  4.095 2.300 4.150 2.640 ;
        RECT  3.390 2.940 4.150 3.260 ;
        RECT  1.535 3.030 3.390 3.260 ;
        RECT  1.455 2.940 1.535 3.260 ;
        RECT  1.440 2.660 1.455 3.260 ;
        RECT  1.100 2.605 1.440 3.260 ;
        RECT  1.085 2.660 1.100 3.260 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 1.680 3.740 2.075 ;
        RECT  2.150 1.745 3.400 2.075 ;
        RECT  1.810 1.745 2.150 2.530 ;
        RECT  1.470 1.745 1.810 2.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.480 2.305 3.200 2.685 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.760 -0.400 7.260 0.400 ;
        RECT  6.420 -0.400 6.760 0.575 ;
        RECT  5.030 -0.400 6.420 0.400 ;
        RECT  4.690 -0.400 5.030 0.575 ;
        RECT  2.000 -0.400 4.690 0.400 ;
        RECT  1.660 -0.400 2.000 0.575 ;
        RECT  0.520 -0.400 1.660 0.400 ;
        RECT  0.180 -0.400 0.520 1.740 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.840 4.640 7.260 5.440 ;
        RECT  6.500 4.465 6.840 5.440 ;
        RECT  5.400 4.640 6.500 5.440 ;
        RECT  5.060 4.465 5.400 5.440 ;
        RECT  0.520 4.640 5.060 5.440 ;
        RECT  0.180 4.040 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.665 2.100 6.720 2.440 ;
        RECT  6.435 0.935 6.665 4.195 ;
        RECT  2.930 0.935 6.435 1.165 ;
        RECT  6.380 2.100 6.435 2.440 ;
        RECT  2.920 3.965 6.435 4.195 ;
        RECT  2.590 0.645 2.930 1.455 ;
        RECT  2.580 3.965 2.920 4.305 ;
        RECT  2.285 0.935 2.590 1.165 ;
        RECT  2.055 0.935 2.285 1.450 ;
        RECT  1.240 1.220 2.055 1.450 ;
        RECT  0.900 0.930 1.240 1.740 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 0.765 3.820 4.240 ;
        RECT  3.390 0.765 3.590 1.575 ;
        RECT  3.430 2.940 3.590 4.240 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.620 2.940 3.160 3.220 ;
        RECT  2.390 2.320 2.620 3.220 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.215 2.000 2.660 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 0.700 1.310 1.110 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.545 2.380 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 -0.400 3.960 0.400 ;
        RECT  1.985 -0.400 2.325 0.575 ;
        RECT  0.520 -0.400 1.985 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.010 4.640 3.960 5.440 ;
        RECT  2.670 4.465 3.010 5.440 ;
        RECT  0.000 4.640 2.670 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.155 1.940 3.305 2.420 ;
        RECT  2.925 1.400 3.155 2.420 ;
        RECT  2.410 1.400 2.925 1.630 ;
        RECT  2.070 1.345 2.410 1.685 ;
        RECT  1.025 1.400 2.070 1.630 ;
        RECT  1.005 1.345 1.025 1.630 ;
        RECT  0.775 1.345 1.005 3.010 ;
        RECT  0.520 2.780 0.775 3.010 ;
        RECT  0.290 2.780 0.520 3.880 ;
        RECT  0.180 3.070 0.290 3.880 ;
    END
END OR4X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.800 3.500 3.820 3.870 ;
        RECT  3.570 0.950 3.800 3.870 ;
        RECT  3.420 0.950 3.570 1.290 ;
        RECT  3.240 3.500 3.570 3.870 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.715 2.330 3.190 2.795 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 2.330 1.980 3.220 ;
        RECT  1.460 2.910 1.750 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.170 1.280 2.665 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.755 0.560 3.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.000 -0.400 3.960 0.400 ;
        RECT  2.660 -0.400 3.000 0.575 ;
        RECT  1.120 -0.400 2.660 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 4.640 3.960 5.440 ;
        RECT  2.480 4.465 2.820 5.440 ;
        RECT  0.000 4.640 2.480 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.480 1.655 3.295 2.005 ;
        RECT  2.250 1.180 2.480 3.915 ;
        RECT  2.060 1.180 2.250 1.520 ;
        RECT  0.540 3.685 2.250 3.915 ;
        RECT  0.800 1.180 2.060 1.410 ;
        RECT  0.570 1.180 0.800 1.780 ;
        RECT  0.460 1.440 0.570 1.780 ;
        RECT  0.200 3.630 0.540 3.970 ;
    END
END OR4X1

MACRO OR3XL
    CLASS CORE ;
    FOREIGN OR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.900 1.460 3.130 3.660 ;
        RECT  2.745 1.460 2.900 1.800 ;
        RECT  2.780 2.965 2.900 3.660 ;
        RECT  2.620 3.320 2.780 3.660 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.675 2.000 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.820 1.475 2.335 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.755 2.670 0.985 4.315 ;
        RECT  0.600 2.670 0.755 3.030 ;
        RECT  0.215 4.085 0.755 4.315 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 -0.400 3.300 0.400 ;
        RECT  2.180 -0.400 2.520 0.575 ;
        RECT  0.560 -0.400 2.180 0.400 ;
        RECT  0.220 -0.400 0.560 0.575 ;
        RECT  0.000 -0.400 0.220 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 4.640 3.300 5.440 ;
        RECT  2.060 4.465 2.400 5.440 ;
        RECT  0.000 4.640 2.060 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.330 2.090 2.670 2.430 ;
        RECT  2.300 2.090 2.330 2.320 ;
        RECT  2.070 1.235 2.300 2.320 ;
        RECT  1.820 1.235 2.070 1.465 ;
        RECT  1.480 0.805 1.820 1.465 ;
        RECT  0.520 1.235 1.480 1.465 ;
        RECT  0.370 1.235 0.520 1.800 ;
        RECT  0.370 3.265 0.520 3.605 ;
        RECT  0.140 1.235 0.370 3.605 ;
    END
END OR3XL

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR3XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 2.850 4.970 3.220 ;
        RECT  4.480 1.390 4.730 1.730 ;
        RECT  4.100 1.390 4.480 3.220 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 1.735 3.585 1.965 ;
        RECT  3.175 1.735 3.405 3.185 ;
        RECT  3.085 2.940 3.175 3.185 ;
        RECT  2.855 2.955 3.085 3.185 ;
        RECT  2.585 2.955 2.855 3.220 ;
        RECT  2.355 2.955 2.585 3.375 ;
        RECT  0.875 3.145 2.355 3.375 ;
        RECT  0.800 2.940 0.875 3.375 ;
        RECT  0.570 2.535 0.800 3.375 ;
        RECT  0.460 2.535 0.570 3.255 ;
        RECT  0.140 2.860 0.460 3.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 1.920 2.815 2.450 ;
        RECT  1.105 1.920 2.475 2.150 ;
        RECT  0.980 1.845 1.105 2.150 ;
        RECT  0.640 1.810 0.980 2.150 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 2.380 2.035 2.915 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.550 -0.400 5.940 0.400 ;
        RECT  5.210 -0.400 5.550 0.575 ;
        RECT  3.895 -0.400 5.210 0.400 ;
        RECT  3.555 -0.400 3.895 0.575 ;
        RECT  2.305 -0.400 3.555 0.400 ;
        RECT  1.965 -0.400 2.305 0.995 ;
        RECT  0.000 -0.400 1.965 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.605 4.640 5.940 5.440 ;
        RECT  5.265 4.065 5.605 5.440 ;
        RECT  4.280 4.640 5.265 5.440 ;
        RECT  3.940 4.065 4.280 5.440 ;
        RECT  0.520 4.640 3.940 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.200 0.895 5.430 3.770 ;
        RECT  3.100 0.895 5.200 1.125 ;
        RECT  4.945 2.235 5.200 2.575 ;
        RECT  3.165 3.540 5.200 3.770 ;
        RECT  2.935 3.540 3.165 3.995 ;
        RECT  3.085 0.895 3.100 1.505 ;
        RECT  2.745 0.680 3.085 1.505 ;
        RECT  2.400 3.765 2.935 3.995 ;
        RECT  1.535 1.275 2.745 1.505 ;
        RECT  2.060 3.765 2.400 4.105 ;
        RECT  1.195 0.680 1.535 1.505 ;
    END
END OR3X4

MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR3XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.740 0.765 3.820 2.100 ;
        RECT  3.510 0.765 3.740 4.240 ;
        RECT  3.440 0.765 3.510 2.100 ;
        RECT  3.400 2.960 3.510 4.240 ;
        RECT  3.400 0.765 3.440 1.575 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 2.525 2.520 3.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.775 1.940 2.130 ;
        RECT  1.480 1.775 1.820 2.175 ;
        RECT  1.380 1.775 1.480 2.130 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 2.380 1.160 2.805 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 -0.400 3.960 0.400 ;
        RECT  2.680 -0.400 3.020 0.950 ;
        RECT  1.350 -0.400 2.680 0.400 ;
        RECT  1.010 -0.400 1.350 0.575 ;
        RECT  0.000 -0.400 1.010 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 4.640 3.960 5.440 ;
        RECT  2.600 4.465 2.940 5.440 ;
        RECT  0.000 4.640 2.600 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.065 2.020 3.105 2.385 ;
        RECT  2.835 1.315 3.065 2.385 ;
        RECT  0.530 1.315 2.835 1.545 ;
        RECT  0.580 3.175 0.920 3.985 ;
        RECT  0.395 3.175 0.580 3.405 ;
        RECT  0.395 1.260 0.530 1.600 ;
        RECT  0.165 1.260 0.395 3.405 ;
    END
END OR3X2

MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR3XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.585 2.330 3.825 2.965 ;
        RECT  3.585 1.060 3.590 1.400 ;
        RECT  3.355 1.060 3.585 3.685 ;
        RECT  3.250 1.060 3.355 1.415 ;
        RECT  3.170 2.875 3.355 3.685 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 2.570 2.500 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.335 1.730 1.840 2.150 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.705 2.380 1.210 2.930 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.700 -0.400 3.960 0.400 ;
        RECT  2.360 -0.400 2.700 0.575 ;
        RECT  1.370 -0.400 2.360 0.400 ;
        RECT  1.030 -0.400 1.370 0.575 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 4.640 3.960 5.440 ;
        RECT  2.355 4.465 2.695 5.440 ;
        RECT  0.000 4.640 2.355 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.930 1.770 3.080 2.110 ;
        RECT  2.630 1.200 2.930 2.110 ;
        RECT  2.000 1.200 2.630 1.500 ;
        RECT  1.660 1.150 2.000 1.500 ;
        RECT  0.540 1.200 1.660 1.500 ;
        RECT  0.395 3.320 0.720 3.685 ;
        RECT  0.395 1.150 0.540 1.500 ;
        RECT  0.165 1.150 0.395 3.685 ;
    END
END OR3X1

MACRO OR2XL
    CLASS CORE ;
    FOREIGN OR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.250 1.430 2.480 3.640 ;
        RECT  2.120 1.430 2.250 1.770 ;
        RECT  2.120 2.920 2.250 3.640 ;
        RECT  2.085 3.300 2.120 3.640 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 2.380 1.220 3.220 ;
        RECT  0.860 2.380 1.180 3.240 ;
        RECT  0.800 2.940 0.860 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.160 1.990 0.580 2.680 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.390 -0.400 2.640 0.400 ;
        RECT  0.450 -0.400 1.390 0.575 ;
        RECT  0.000 -0.400 0.450 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.450 4.640 2.640 5.440 ;
        RECT  1.110 4.410 1.450 5.440 ;
        RECT  0.000 4.640 1.110 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.775 2.150 2.020 2.490 ;
        RECT  1.545 1.315 1.775 3.805 ;
        RECT  0.810 1.315 1.545 1.545 ;
        RECT  0.540 3.575 1.545 3.805 ;
        RECT  0.445 1.315 0.810 1.700 ;
        RECT  0.200 3.520 0.540 3.860 ;
    END
END OR2XL

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR2XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 1.360 2.640 1.700 ;
        RECT  2.505 2.740 2.520 3.080 ;
        RECT  2.500 2.620 2.505 3.080 ;
        RECT  2.180 1.260 2.500 3.080 ;
        RECT  2.120 1.260 2.180 2.660 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 2.010 1.840 2.785 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.645 0.520 2.335 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 -0.400 3.960 0.400 ;
        RECT  2.980 -0.400 3.320 0.575 ;
        RECT  2.000 -0.400 2.980 0.400 ;
        RECT  1.660 -0.400 2.000 0.960 ;
        RECT  0.520 -0.400 1.660 0.400 ;
        RECT  0.180 -0.400 0.520 1.280 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 4.640 3.960 5.440 ;
        RECT  2.860 4.465 3.200 5.440 ;
        RECT  1.840 4.640 2.860 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.010 2.100 3.120 2.440 ;
        RECT  2.780 2.100 3.010 3.540 ;
        RECT  1.000 3.310 2.780 3.540 ;
        RECT  1.000 1.160 1.240 1.500 ;
        RECT  0.770 1.160 1.000 3.540 ;
        RECT  0.180 2.810 0.770 3.150 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR2XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.220 0.825 2.450 3.840 ;
        RECT  2.065 0.825 2.220 1.635 ;
        RECT  2.060 3.030 2.220 3.840 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.740 1.270 2.345 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.650 0.520 2.285 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 2.640 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 4.640 2.640 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.000 4.640 1.300 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.735 2.110 1.990 2.450 ;
        RECT  1.505 1.170 1.735 3.260 ;
        RECT  1.080 1.170 1.505 1.400 ;
        RECT  0.520 3.030 1.505 3.260 ;
        RECT  0.740 1.060 1.080 1.400 ;
        RECT  0.180 3.030 0.520 3.370 ;
    END
END OR2X2

MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR2XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.250 1.320 2.480 3.640 ;
        RECT  2.120 1.320 2.250 1.660 ;
        RECT  2.120 2.920 2.250 3.640 ;
        RECT  2.085 3.300 2.120 3.640 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 2.380 1.220 3.220 ;
        RECT  0.860 2.380 1.180 3.240 ;
        RECT  0.800 2.940 0.860 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.160 1.990 0.580 2.680 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.390 -0.400 2.640 0.400 ;
        RECT  0.450 -0.400 1.390 0.575 ;
        RECT  0.000 -0.400 0.450 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.450 4.640 2.640 5.440 ;
        RECT  1.095 4.385 1.450 5.440 ;
        RECT  0.000 4.640 1.095 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.775 2.150 2.020 2.490 ;
        RECT  1.545 1.315 1.775 3.805 ;
        RECT  0.810 1.315 1.545 1.545 ;
        RECT  0.540 3.575 1.545 3.805 ;
        RECT  0.445 1.315 0.810 1.700 ;
        RECT  0.200 3.520 0.540 3.860 ;
    END
END OR2X1

MACRO OAI33XL
    CLASS CORE ;
    FOREIGN OAI33XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.255 5.065 3.725 ;
        RECT  4.465 1.255 4.835 1.485 ;
        RECT  2.020 3.495 4.835 3.725 ;
        RECT  4.235 1.255 4.465 1.805 ;
        RECT  3.185 1.575 4.235 1.805 ;
        RECT  2.955 1.200 3.185 1.805 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.520 3.050 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.085 1.265 2.660 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 2.505 1.935 3.195 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.050 2.100 4.480 2.635 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.060 2.210 3.745 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.605 2.940 3.085 3.195 ;
        RECT  2.375 2.625 2.605 3.195 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 -0.400 5.280 0.400 ;
        RECT  1.460 -0.400 1.800 1.345 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.240 4.640 5.280 5.440 ;
        RECT  3.900 4.465 4.240 5.440 ;
        RECT  0.520 4.640 3.900 5.440 ;
        RECT  0.180 3.485 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.825 1.115 3.960 1.345 ;
        RECT  3.595 0.735 3.825 1.345 ;
        RECT  2.465 0.735 3.595 0.965 ;
        RECT  2.235 0.735 2.465 1.810 ;
        RECT  1.025 1.580 2.235 1.810 ;
        RECT  0.795 1.170 1.025 1.810 ;
    END
END OAI33XL

MACRO OAI33X4
    CLASS CORE ;
    FOREIGN OAI33X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI33XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.650 1.820 5.800 3.220 ;
        RECT  5.420 1.420 5.650 3.220 ;
        RECT  5.065 1.420 5.420 1.650 ;
        RECT  4.715 2.795 5.420 3.025 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 2.600 4.405 3.195 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 1.780 3.820 2.135 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.315 2.405 3.085 2.940 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.530 2.360 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.405 1.375 2.940 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 3.920 2.160 4.405 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.085 -0.400 7.260 0.400 ;
        RECT  5.745 -0.400 6.085 0.575 ;
        RECT  4.725 -0.400 5.745 0.400 ;
        RECT  4.385 -0.400 4.725 0.575 ;
        RECT  3.165 -0.400 4.385 0.400 ;
        RECT  2.825 -0.400 3.165 0.575 ;
        RECT  0.000 -0.400 2.825 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.695 4.640 7.260 5.440 ;
        RECT  5.355 4.090 5.695 5.440 ;
        RECT  4.305 4.640 5.355 5.440 ;
        RECT  3.965 4.465 4.305 5.440 ;
        RECT  0.520 4.640 3.965 5.440 ;
        RECT  0.180 3.420 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.725 1.365 6.850 1.705 ;
        RECT  6.495 0.885 6.725 3.410 ;
        RECT  4.760 0.885 6.495 1.115 ;
        RECT  6.035 2.540 6.265 3.715 ;
        RECT  3.435 3.485 6.035 3.715 ;
        RECT  4.530 0.885 4.760 2.235 ;
        RECT  2.220 1.235 3.880 1.465 ;
        RECT  3.205 3.275 3.435 3.715 ;
        RECT  1.845 3.275 3.205 3.505 ;
        RECT  1.615 1.235 1.845 3.505 ;
        RECT  0.180 1.235 1.615 1.465 ;
    END
END OAI33X4

MACRO OAI33X2
    CLASS CORE ;
    FOREIGN OAI33X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI33XL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.895 1.360 8.125 3.755 ;
        RECT  4.715 1.360 7.895 1.590 ;
        RECT  7.705 3.500 7.895 3.755 ;
        RECT  6.120 3.525 7.705 3.755 ;
        RECT  5.780 3.525 6.120 4.410 ;
        RECT  2.360 3.525 5.780 3.755 ;
        RECT  2.020 3.470 2.360 3.810 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.830 2.245 3.940 2.585 ;
        RECT  3.600 2.245 3.830 3.140 ;
        RECT  0.520 2.910 3.600 3.140 ;
        RECT  0.520 2.250 0.530 2.590 ;
        RECT  0.290 2.250 0.520 3.140 ;
        RECT  0.215 2.250 0.290 2.635 ;
        RECT  0.190 2.250 0.215 2.590 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.215 1.820 3.270 2.335 ;
        RECT  2.855 1.820 3.215 2.635 ;
        RECT  1.430 1.820 2.855 2.050 ;
        RECT  1.095 1.820 1.430 2.335 ;
        RECT  1.090 1.995 1.095 2.335 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 2.305 2.500 2.660 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.435 2.380 7.665 3.195 ;
        RECT  4.405 2.965 7.435 3.195 ;
        RECT  4.405 1.260 4.410 1.910 ;
        RECT  4.175 1.260 4.405 3.195 ;
        RECT  4.070 1.260 4.175 1.910 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.635 1.920 6.865 2.330 ;
        RECT  5.065 1.920 6.635 2.150 ;
        RECT  5.025 1.845 5.065 2.150 ;
        RECT  4.795 1.845 5.025 2.330 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 2.380 6.190 2.735 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 -0.400 8.580 0.400 ;
        RECT  2.030 -0.400 2.370 0.950 ;
        RECT  0.520 -0.400 2.030 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.000 4.640 8.580 5.440 ;
        RECT  7.660 4.465 8.000 5.440 ;
        RECT  4.240 4.640 7.660 5.440 ;
        RECT  3.900 4.465 4.240 5.440 ;
        RECT  0.520 4.640 3.900 5.440 ;
        RECT  0.180 3.370 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.370 0.665 7.795 0.895 ;
        RECT  3.140 0.665 3.370 1.590 ;
        RECT  0.970 1.360 3.140 1.590 ;
    END
END OAI33X2

MACRO OAI33X1
    CLASS CORE ;
    FOREIGN OAI33X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI33XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.940 2.405 5.065 2.635 ;
        RECT  4.710 1.125 4.940 3.725 ;
        RECT  4.500 1.125 4.710 1.740 ;
        RECT  2.360 3.495 4.710 3.725 ;
        RECT  3.400 1.510 4.500 1.740 ;
        RECT  3.060 1.315 3.400 1.740 ;
        RECT  2.020 3.440 2.360 3.780 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.950 0.530 2.660 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.970 1.430 2.660 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 2.255 2.150 2.595 ;
        RECT  1.810 2.255 2.040 3.195 ;
        RECT  1.535 2.940 1.810 3.195 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 2.965 4.405 3.195 ;
        RECT  4.335 2.185 4.390 2.525 ;
        RECT  4.105 2.185 4.335 3.195 ;
        RECT  4.050 2.185 4.105 2.525 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.260 2.120 3.820 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 2.965 3.085 3.195 ;
        RECT  2.720 2.250 2.950 3.195 ;
        RECT  2.535 2.250 2.720 2.590 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 -0.400 5.280 0.400 ;
        RECT  1.620 -0.400 1.960 1.275 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 1.450 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.590 4.640 5.280 5.440 ;
        RECT  4.250 4.465 4.590 5.440 ;
        RECT  0.520 4.640 4.250 5.440 ;
        RECT  0.180 3.295 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 0.845 4.120 1.275 ;
        RECT  2.680 0.845 3.780 1.075 ;
        RECT  2.570 0.845 2.680 1.470 ;
        RECT  2.450 0.845 2.570 1.735 ;
        RECT  2.340 1.130 2.450 1.735 ;
        RECT  1.240 1.505 2.340 1.735 ;
        RECT  1.010 1.105 1.240 1.735 ;
        RECT  0.900 1.105 1.010 1.445 ;
    END
END OAI33X1

MACRO OAI32XL
    CLASS CORE ;
    FOREIGN OAI32XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.675 4.405 3.890 ;
        RECT  3.545 1.675 4.175 1.905 ;
        RECT  2.360 3.660 4.175 3.890 ;
        RECT  3.315 1.130 3.545 1.905 ;
        RECT  3.060 1.130 3.315 1.360 ;
        RECT  2.020 3.605 2.360 3.945 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 2.380 3.820 3.145 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 2.180 3.160 2.660 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.265 0.530 2.995 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 1.995 1.480 2.335 ;
        RECT  0.800 1.995 1.275 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 2.665 2.120 3.220 ;
        RECT  1.460 2.940 1.655 3.220 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 -0.400 4.620 0.400 ;
        RECT  1.620 -0.400 1.960 1.275 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 1.275 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.680 4.640 4.620 5.440 ;
        RECT  3.340 4.465 3.680 5.440 ;
        RECT  0.520 4.640 3.340 5.440 ;
        RECT  0.180 3.295 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.010 0.935 4.120 1.275 ;
        RECT  3.780 0.630 4.010 1.275 ;
        RECT  2.680 0.630 3.780 0.860 ;
        RECT  2.570 0.630 2.680 1.415 ;
        RECT  2.450 0.630 2.570 1.765 ;
        RECT  2.340 1.075 2.450 1.765 ;
        RECT  1.240 1.535 2.340 1.765 ;
        RECT  1.010 1.075 1.240 1.765 ;
        RECT  0.900 1.075 1.010 1.415 ;
    END
END OAI32XL

MACRO OAI32X4
    CLASS CORE ;
    FOREIGN OAI32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI32XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.990 1.820 5.140 3.220 ;
        RECT  4.760 1.460 4.990 3.220 ;
        RECT  4.440 1.460 4.760 1.690 ;
        RECT  4.175 2.890 4.760 3.120 ;
        RECT  4.100 1.350 4.440 1.690 ;
        RECT  3.825 2.890 4.175 3.230 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.520 3.110 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 4.010 1.435 4.405 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 2.380 3.820 2.660 ;
        RECT  2.900 2.210 3.240 2.660 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 2.965 3.085 3.195 ;
        RECT  2.320 2.215 2.550 3.195 ;
        RECT  2.210 2.215 2.320 2.555 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 2.380 1.840 3.010 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.120 -0.400 6.600 0.400 ;
        RECT  4.780 -0.400 5.120 0.575 ;
        RECT  3.690 -0.400 4.780 0.400 ;
        RECT  3.350 -0.400 3.690 0.575 ;
        RECT  2.560 -0.400 3.350 0.400 ;
        RECT  2.220 -0.400 2.560 0.575 ;
        RECT  0.000 -0.400 2.220 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.980 4.640 6.600 5.440 ;
        RECT  4.640 4.090 4.980 5.440 ;
        RECT  3.525 4.640 4.640 5.440 ;
        RECT  3.185 4.090 3.525 5.440 ;
        RECT  0.520 4.640 3.185 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.835 0.815 6.065 3.410 ;
        RECT  5.545 0.815 5.835 1.275 ;
        RECT  5.370 2.540 5.600 3.695 ;
        RECT  3.810 0.815 5.545 1.045 ;
        RECT  1.640 3.465 5.370 3.695 ;
        RECT  4.050 1.920 4.390 2.260 ;
        RECT  3.810 1.920 4.050 2.150 ;
        RECT  3.580 0.815 3.810 2.150 ;
        RECT  2.780 1.260 3.120 1.600 ;
        RECT  1.800 1.315 2.780 1.545 ;
        RECT  1.460 1.260 1.800 1.600 ;
        RECT  1.300 3.395 1.640 3.735 ;
        RECT  0.980 3.395 1.300 3.625 ;
        RECT  0.980 1.260 1.080 1.600 ;
        RECT  0.750 1.260 0.980 3.625 ;
        RECT  0.740 1.260 0.750 1.600 ;
    END
END OAI32X4

MACRO OAI32X2
    CLASS CORE ;
    FOREIGN OAI32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI32XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.385 1.495 6.615 4.050 ;
        RECT  6.155 1.495 6.385 1.725 ;
        RECT  6.080 3.525 6.385 4.050 ;
        RECT  5.900 1.440 6.155 1.725 ;
        RECT  5.565 3.820 6.080 4.050 ;
        RECT  5.560 1.440 5.900 1.780 ;
        RECT  5.225 3.765 5.565 4.105 ;
        RECT  4.250 1.495 5.560 1.725 ;
        RECT  3.570 3.820 5.225 4.050 ;
        RECT  3.910 1.440 4.250 1.780 ;
        RECT  3.340 3.820 3.570 4.355 ;
        RECT  3.085 4.060 3.340 4.355 ;
        RECT  2.360 4.125 3.085 4.355 ;
        RECT  2.020 4.070 2.360 4.410 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.655 2.010 5.995 2.350 ;
        RECT  4.520 2.010 5.655 2.240 ;
        RECT  4.405 2.010 4.520 2.615 ;
        RECT  4.175 2.010 4.405 2.635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.800 2.510 5.325 3.195 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 2.580 3.830 2.965 ;
        RECT  3.490 2.580 3.720 3.240 ;
        RECT  2.815 3.010 3.490 3.240 ;
        RECT  2.585 3.010 2.815 3.725 ;
        RECT  1.225 3.495 2.585 3.725 ;
        RECT  0.995 2.685 1.225 3.725 ;
        RECT  0.760 2.685 0.995 2.965 ;
        RECT  0.705 2.575 0.760 2.965 ;
        RECT  0.420 2.405 0.705 2.965 ;
        RECT  0.215 2.405 0.420 2.635 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 2.010 3.160 2.650 ;
        RECT  2.780 2.065 2.820 2.650 ;
        RECT  1.435 2.065 2.780 2.295 ;
        RECT  1.095 2.010 1.435 2.350 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 2.580 2.120 3.195 ;
        RECT  1.535 2.965 1.680 3.195 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.530 -0.400 7.260 0.400 ;
        RECT  2.190 -0.400 2.530 0.950 ;
        RECT  0.680 -0.400 2.190 0.400 ;
        RECT  0.340 -0.400 0.680 0.950 ;
        RECT  0.000 -0.400 0.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.885 4.640 7.260 5.440 ;
        RECT  6.545 4.465 6.885 5.440 ;
        RECT  4.245 4.640 6.545 5.440 ;
        RECT  3.905 4.465 4.245 5.440 ;
        RECT  0.520 4.640 3.905 5.440 ;
        RECT  0.180 3.620 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.455 0.630 5.265 0.970 ;
        RECT  3.380 0.685 4.455 0.915 ;
        RECT  3.150 0.685 3.380 1.780 ;
        RECT  3.040 1.440 3.150 1.780 ;
        RECT  1.790 1.495 3.040 1.725 ;
        RECT  0.980 1.440 1.790 1.780 ;
    END
END OAI32X2

MACRO OAI32X1
    CLASS CORE ;
    FOREIGN OAI32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI32XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.510 4.405 3.680 ;
        RECT  4.100 1.510 4.175 1.845 ;
        RECT  2.020 3.450 4.175 3.680 ;
        RECT  3.400 1.510 4.100 1.740 ;
        RECT  3.060 1.320 3.400 1.740 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 2.045 3.820 2.690 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.840 2.965 3.085 3.195 ;
        RECT  2.610 2.275 2.840 3.195 ;
        RECT  2.500 2.275 2.610 2.615 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.530 2.985 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.915 1.430 2.145 ;
        RECT  0.875 1.915 1.180 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 2.575 1.990 3.195 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 -0.400 4.620 0.400 ;
        RECT  1.620 -0.400 1.960 1.225 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 1.280 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.680 4.640 4.620 5.440 ;
        RECT  3.340 4.410 3.680 5.440 ;
        RECT  0.520 4.640 3.340 5.440 ;
        RECT  0.180 4.145 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 0.860 4.120 1.280 ;
        RECT  2.680 0.860 3.780 1.090 ;
        RECT  2.570 0.860 2.680 1.450 ;
        RECT  2.450 0.860 2.570 1.685 ;
        RECT  2.340 1.110 2.450 1.685 ;
        RECT  1.240 1.455 2.340 1.685 ;
        RECT  1.010 1.080 1.240 1.685 ;
        RECT  0.900 1.080 1.010 1.420 ;
    END
END OAI32X1

MACRO OAI31XL
    CLASS CORE ;
    FOREIGN OAI31XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.255 3.745 3.400 ;
        RECT  2.780 1.255 3.515 1.485 ;
        RECT  1.860 3.170 3.515 3.400 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.590 2.380 3.160 2.890 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.530 3.070 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.710 1.705 1.325 2.120 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.735 2.105 2.635 ;
        RECT  1.535 2.405 1.840 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 3.960 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 4.640 3.960 5.440 ;
        RECT  2.620 4.465 2.960 5.440 ;
        RECT  0.520 4.640 2.620 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.740 1.245 2.400 1.475 ;
    END
END OAI31XL

MACRO OAI31X4
    CLASS CORE ;
    FOREIGN OAI31X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI31XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 1.820 4.480 3.220 ;
        RECT  4.100 1.440 4.330 3.220 ;
        RECT  3.880 1.440 4.100 1.670 ;
        RECT  3.640 2.990 4.100 3.220 ;
        RECT  3.540 1.330 3.880 1.670 ;
        RECT  3.410 2.740 3.640 3.220 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 2.240 0.520 2.915 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.995 2.965 3.085 3.195 ;
        RECT  2.765 2.765 2.995 3.195 ;
        RECT  2.600 2.765 2.765 2.995 ;
        RECT  2.260 2.655 2.600 2.995 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 1.675 2.500 2.100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.405 1.765 2.635 ;
        RECT  1.210 1.895 1.505 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.560 -0.400 5.940 0.400 ;
        RECT  4.220 -0.400 4.560 0.575 ;
        RECT  3.200 -0.400 4.220 0.400 ;
        RECT  2.860 -0.400 3.200 0.575 ;
        RECT  1.900 -0.400 2.860 0.400 ;
        RECT  1.560 -0.400 1.900 0.575 ;
        RECT  0.000 -0.400 1.560 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 4.640 5.940 5.440 ;
        RECT  4.000 4.090 4.340 5.440 ;
        RECT  3.055 4.640 4.000 5.440 ;
        RECT  2.715 4.090 3.055 5.440 ;
        RECT  0.520 4.640 2.715 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.180 0.830 5.410 4.225 ;
        RECT  4.980 0.830 5.180 1.170 ;
        RECT  5.065 3.995 5.180 4.225 ;
        RECT  4.725 3.995 5.065 4.335 ;
        RECT  3.175 0.830 4.980 1.060 ;
        RECT  4.720 2.535 4.950 3.680 ;
        RECT  1.090 3.450 4.720 3.680 ;
        RECT  3.300 2.000 3.640 2.340 ;
        RECT  3.175 2.000 3.300 2.230 ;
        RECT  2.945 0.830 3.175 2.230 ;
        RECT  2.220 1.060 2.560 1.400 ;
        RECT  1.240 1.060 2.220 1.290 ;
        RECT  0.900 1.060 1.240 1.400 ;
        RECT  0.980 3.220 1.090 3.680 ;
        RECT  0.750 1.710 0.980 3.680 ;
        RECT  0.520 1.710 0.750 1.940 ;
        RECT  0.290 1.140 0.520 1.940 ;
        RECT  0.180 1.140 0.290 1.480 ;
    END
END OAI31X4

MACRO OAI31X2
    CLASS CORE ;
    FOREIGN OAI31X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI31XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.970 1.440 5.080 1.845 ;
        RECT  4.515 3.375 4.985 3.825 ;
        RECT  4.740 1.440 4.970 2.150 ;
        RECT  4.515 1.920 4.740 2.150 ;
        RECT  4.285 1.920 4.515 3.825 ;
        RECT  4.175 3.525 4.285 3.825 ;
        RECT  2.360 3.595 4.175 3.825 ;
        RECT  2.020 3.595 2.360 4.405 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.760 2.380 5.195 3.020 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.850 2.580 4.020 2.920 ;
        RECT  3.680 2.580 3.850 3.325 ;
        RECT  3.620 2.635 3.680 3.325 ;
        RECT  3.515 2.965 3.620 3.325 ;
        RECT  0.875 3.095 3.515 3.325 ;
        RECT  0.760 2.940 0.875 3.325 ;
        RECT  0.530 2.580 0.760 3.325 ;
        RECT  0.420 2.580 0.530 2.920 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 2.265 3.350 2.605 ;
        RECT  3.010 1.870 3.240 2.605 ;
        RECT  1.765 1.870 3.010 2.100 ;
        RECT  1.535 1.845 1.765 2.100 ;
        RECT  1.460 1.870 1.535 2.100 ;
        RECT  1.230 1.870 1.460 2.605 ;
        RECT  1.090 2.265 1.230 2.605 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 2.380 2.500 2.805 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.800 -0.400 5.940 0.400 ;
        RECT  3.460 -0.400 3.800 0.575 ;
        RECT  2.400 -0.400 3.460 0.400 ;
        RECT  2.060 -0.400 2.400 0.575 ;
        RECT  1.080 -0.400 2.060 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.705 4.640 5.940 5.440 ;
        RECT  5.365 3.385 5.705 5.440 ;
        RECT  4.300 4.640 5.365 5.440 ;
        RECT  3.960 4.465 4.300 5.440 ;
        RECT  0.520 4.640 3.960 5.440 ;
        RECT  0.180 3.620 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 1.410 4.360 1.640 ;
        RECT  2.960 0.635 3.190 1.640 ;
        RECT  2.640 0.635 2.960 1.535 ;
        RECT  1.840 1.305 2.640 1.535 ;
        RECT  1.500 1.250 1.840 1.590 ;
        RECT  0.520 1.360 1.500 1.590 ;
        RECT  0.180 1.250 0.520 1.590 ;
    END
END OAI31X2

MACRO OAI31X1
    CLASS CORE ;
    FOREIGN OAI31X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI31XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 0.990 3.745 3.550 ;
        RECT  3.440 0.990 3.515 1.285 ;
        RECT  3.440 3.195 3.515 3.550 ;
        RECT  3.140 0.990 3.440 1.220 ;
        RECT  2.060 3.320 3.440 3.550 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.850 3.185 2.635 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.020 0.520 2.660 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.820 1.480 2.130 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 2.305 2.170 2.735 ;
        RECT  1.535 2.395 1.750 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 -0.400 3.960 0.400 ;
        RECT  2.000 -0.400 2.040 0.430 ;
        RECT  1.660 -0.400 2.000 0.575 ;
        RECT  1.620 -0.400 1.660 0.430 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 4.640 3.960 5.440 ;
        RECT  2.620 4.465 2.960 5.440 ;
        RECT  0.520 4.640 2.620 5.440 ;
        RECT  0.180 3.820 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.900 1.245 2.760 1.475 ;
    END
END OAI31X1

MACRO OAI2BB2XL
    CLASS CORE ;
    FOREIGN OAI2BB2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 1.845 4.405 2.075 ;
        RECT  4.150 0.930 4.380 3.580 ;
        RECT  4.040 0.930 4.150 1.270 ;
        RECT  4.100 3.195 4.150 3.580 ;
        RECT  2.880 3.350 4.100 3.580 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.025 2.160 2.500 2.660 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.730 1.820 3.160 2.500 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.985 2.090 1.215 2.660 ;
        RECT  0.830 2.100 0.985 2.660 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.645 0.600 2.130 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 -0.400 4.620 0.400 ;
        RECT  2.600 -0.400 2.940 1.075 ;
        RECT  0.520 -0.400 2.600 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 4.640 4.620 5.440 ;
        RECT  3.640 4.465 3.980 5.440 ;
        RECT  2.000 4.640 3.640 5.440 ;
        RECT  1.660 4.465 2.000 5.440 ;
        RECT  0.700 4.640 1.660 5.440 ;
        RECT  0.645 4.465 0.700 5.440 ;
        RECT  0.415 4.410 0.645 5.440 ;
        RECT  0.360 4.465 0.415 5.440 ;
        RECT  0.000 4.640 0.360 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.615 1.840 3.845 3.120 ;
        RECT  3.550 0.790 3.660 1.130 ;
        RECT  1.675 2.890 3.615 3.120 ;
        RECT  3.320 0.790 3.550 1.535 ;
        RECT  2.180 1.305 3.320 1.535 ;
        RECT  1.950 0.655 2.180 1.535 ;
        RECT  1.840 0.655 1.950 0.885 ;
        RECT  1.675 1.300 1.680 1.640 ;
        RECT  1.445 1.300 1.675 3.280 ;
        RECT  1.340 1.300 1.445 1.640 ;
        RECT  1.300 3.050 1.445 3.280 ;
        RECT  0.960 3.050 1.300 3.390 ;
    END
END OAI2BB2XL

MACRO OAI2BB2X4
    CLASS CORE ;
    FOREIGN OAI2BB2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB2XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.610 1.170 9.720 1.510 ;
        RECT  9.380 0.805 9.610 2.065 ;
        RECT  5.635 0.805 9.380 1.035 ;
        RECT  9.100 1.835 9.380 2.065 ;
        RECT  8.720 1.820 9.100 3.470 ;
        RECT  6.170 3.130 8.720 3.470 ;
        RECT  5.935 2.945 6.170 3.470 ;
        RECT  4.475 2.945 5.935 3.175 ;
        RECT  5.295 0.660 5.635 1.035 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 2.375 7.265 2.605 ;
        RECT  6.970 2.375 7.045 2.640 ;
        RECT  6.815 2.375 6.970 2.715 ;
        RECT  6.740 2.410 6.815 2.715 ;
        RECT  3.795 2.485 6.740 2.715 ;
        RECT  3.455 2.240 3.795 2.715 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.365 1.915 8.490 2.405 ;
        RECT  8.135 1.915 8.365 2.635 ;
        RECT  6.510 1.915 8.135 2.145 ;
        RECT  6.450 1.915 6.510 2.225 ;
        RECT  6.275 1.915 6.450 2.255 ;
        RECT  6.165 1.995 6.275 2.255 ;
        RECT  4.235 2.025 6.165 2.255 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 2.330 1.630 2.670 ;
        RECT  1.100 2.330 1.290 2.660 ;
        RECT  0.825 2.380 1.100 2.660 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 1.865 2.840 2.205 ;
        RECT  2.500 0.775 2.555 2.205 ;
        RECT  2.325 0.775 2.500 2.095 ;
        RECT  1.155 0.775 2.325 1.005 ;
        RECT  0.925 0.775 1.155 2.020 ;
        RECT  0.875 1.790 0.925 2.020 ;
        RECT  0.610 1.790 0.875 2.100 ;
        RECT  0.270 1.790 0.610 2.130 ;
        RECT  0.215 1.845 0.270 2.075 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.320 -0.400 9.900 0.400 ;
        RECT  7.980 -0.400 8.320 0.575 ;
        RECT  6.955 -0.400 7.980 0.400 ;
        RECT  6.615 -0.400 6.955 0.575 ;
        RECT  4.235 -0.400 6.615 0.400 ;
        RECT  2.785 -0.400 4.235 0.575 ;
        RECT  0.520 -0.400 2.785 0.400 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.680 4.640 9.900 5.440 ;
        RECT  9.340 4.465 9.680 5.440 ;
        RECT  7.595 4.640 9.340 5.440 ;
        RECT  7.255 4.465 7.595 5.440 ;
        RECT  5.515 4.640 7.255 5.440 ;
        RECT  5.175 4.465 5.515 5.440 ;
        RECT  3.495 4.640 5.175 5.440 ;
        RECT  3.155 4.465 3.495 5.440 ;
        RECT  1.990 4.640 3.155 5.440 ;
        RECT  1.650 4.465 1.990 5.440 ;
        RECT  0.520 4.640 1.650 5.440 ;
        RECT  0.180 3.260 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.330 2.295 9.670 4.225 ;
        RECT  5.640 3.885 9.330 4.225 ;
        RECT  8.355 1.360 9.000 1.590 ;
        RECT  8.125 1.360 8.355 1.685 ;
        RECT  4.995 1.455 8.125 1.685 ;
        RECT  5.300 3.420 5.640 4.225 ;
        RECT  4.225 3.420 5.300 3.760 ;
        RECT  4.655 1.390 4.995 1.730 ;
        RECT  3.660 1.455 4.655 1.685 ;
        RECT  3.885 3.090 4.225 3.760 ;
        RECT  2.090 3.090 3.885 3.430 ;
        RECT  3.320 1.390 3.660 1.730 ;
        RECT  1.860 1.345 2.090 3.430 ;
        RECT  1.800 1.345 1.860 1.575 ;
        RECT  0.900 3.090 1.860 3.430 ;
        RECT  1.460 1.235 1.800 1.575 ;
    END
END OAI2BB2X4

MACRO OAI2BB2X2
    CLASS CORE ;
    FOREIGN OAI2BB2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB2XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.155 1.705 6.385 3.875 ;
        RECT  4.515 1.705 6.155 1.935 ;
        RECT  4.825 3.645 6.155 3.875 ;
        RECT  4.485 3.645 4.825 3.985 ;
        RECT  4.285 1.265 4.515 1.935 ;
        RECT  3.305 3.645 4.485 3.875 ;
        RECT  4.040 1.265 4.285 1.495 ;
        RECT  2.965 3.645 3.305 3.985 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.650 2.630 5.805 3.195 ;
        RECT  5.575 2.630 5.650 3.365 ;
        RECT  5.420 2.965 5.575 3.365 ;
        RECT  4.545 3.135 5.420 3.365 ;
        RECT  4.315 2.655 4.545 3.365 ;
        RECT  4.100 2.655 4.315 2.965 ;
        RECT  2.380 2.655 4.100 2.885 ;
        RECT  2.150 2.220 2.380 2.885 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.025 2.675 5.190 2.905 ;
        RECT  4.795 2.185 5.025 2.905 ;
        RECT  3.375 2.185 4.795 2.415 ;
        RECT  3.145 1.845 3.375 2.415 ;
        RECT  2.855 1.845 3.145 2.075 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.460 2.900 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.630 0.760 2.150 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.660 -0.400 6.600 0.400 ;
        RECT  5.320 -0.400 5.660 0.575 ;
        RECT  2.900 -0.400 5.320 0.400 ;
        RECT  2.560 -0.400 2.900 0.575 ;
        RECT  0.520 -0.400 2.560 0.400 ;
        RECT  0.180 -0.400 0.520 1.275 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.145 4.640 6.600 5.440 ;
        RECT  5.805 4.465 6.145 5.440 ;
        RECT  4.065 4.640 5.805 5.440 ;
        RECT  3.725 4.465 4.065 5.440 ;
        RECT  2.025 4.640 3.725 5.440 ;
        RECT  1.685 3.725 2.025 5.440 ;
        RECT  0.585 4.640 1.685 5.440 ;
        RECT  0.245 3.430 0.585 5.440 ;
        RECT  0.000 4.640 0.245 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.080 0.945 6.420 1.285 ;
        RECT  5.100 1.055 6.080 1.285 ;
        RECT  4.985 1.055 5.100 1.475 ;
        RECT  4.755 0.775 4.985 1.475 ;
        RECT  3.660 0.775 4.755 1.005 ;
        RECT  1.920 3.115 3.680 3.345 ;
        RECT  3.320 0.775 3.660 1.115 ;
        RECT  2.545 0.885 3.320 1.115 ;
        RECT  2.315 0.885 2.545 1.585 ;
        RECT  2.000 1.355 2.315 1.585 ;
        RECT  1.770 1.885 1.920 3.495 ;
        RECT  1.770 0.655 1.840 0.885 ;
        RECT  1.690 0.655 1.770 3.495 ;
        RECT  1.435 0.655 1.690 2.115 ;
        RECT  1.305 3.265 1.690 3.495 ;
        RECT  0.965 3.265 1.305 3.630 ;
    END
END OAI2BB2X2

MACRO OAI2BB2X1
    CLASS CORE ;
    FOREIGN OAI2BB2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 1.845 4.405 2.075 ;
        RECT  4.150 1.050 4.380 3.580 ;
        RECT  4.040 1.050 4.150 1.390 ;
        RECT  4.100 3.195 4.150 3.580 ;
        RECT  2.880 3.350 4.100 3.580 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.025 2.160 2.500 2.660 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.730 1.820 3.160 2.500 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.830 2.100 1.215 2.660 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.645 0.600 2.130 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 -0.400 4.620 0.400 ;
        RECT  2.600 -0.400 2.940 0.955 ;
        RECT  0.520 -0.400 2.600 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 4.640 4.620 5.440 ;
        RECT  3.640 4.465 3.980 5.440 ;
        RECT  2.000 4.640 3.640 5.440 ;
        RECT  1.660 4.465 2.000 5.440 ;
        RECT  0.700 4.640 1.660 5.440 ;
        RECT  0.645 4.465 0.700 5.440 ;
        RECT  0.415 4.410 0.645 5.440 ;
        RECT  0.360 4.465 0.415 5.440 ;
        RECT  0.000 4.640 0.360 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.615 1.840 3.845 3.120 ;
        RECT  3.550 0.790 3.660 1.130 ;
        RECT  1.675 2.890 3.615 3.120 ;
        RECT  3.320 0.790 3.550 1.415 ;
        RECT  2.180 1.185 3.320 1.415 ;
        RECT  1.950 0.655 2.180 1.415 ;
        RECT  1.840 0.655 1.950 0.885 ;
        RECT  1.675 1.300 1.680 1.640 ;
        RECT  1.445 1.300 1.675 3.280 ;
        RECT  1.340 1.300 1.445 1.640 ;
        RECT  1.300 3.050 1.445 3.280 ;
        RECT  0.960 3.050 1.300 3.390 ;
    END
END OAI2BB2X1

MACRO OAI2BB1XL
    CLASS CORE ;
    FOREIGN OAI2BB1XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.440 3.155 3.755 ;
        RECT  2.780 1.440 2.925 1.780 ;
        RECT  2.855 3.475 2.925 3.755 ;
        RECT  2.485 3.475 2.855 3.705 ;
        RECT  2.145 3.475 2.485 3.815 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.385 2.380 2.075 2.780 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.485 0.520 3.225 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 1.630 1.180 2.100 ;
        RECT  0.615 1.630 0.955 2.235 ;
        RECT  0.610 1.630 0.615 2.100 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.880 -0.400 3.300 0.400 ;
        RECT  1.540 -0.400 1.880 0.575 ;
        RECT  0.000 -0.400 1.540 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.045 4.640 3.300 5.440 ;
        RECT  2.990 4.465 3.045 5.440 ;
        RECT  2.760 4.410 2.990 5.440 ;
        RECT  2.705 4.465 2.760 5.440 ;
        RECT  1.720 4.640 2.705 5.440 ;
        RECT  0.180 4.465 1.720 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.550 2.100 2.695 2.450 ;
        RECT  2.320 0.985 2.550 3.240 ;
        RECT  0.520 0.985 2.320 1.215 ;
        RECT  1.120 3.010 2.320 3.240 ;
        RECT  0.890 3.010 1.120 3.540 ;
        RECT  0.780 3.200 0.890 3.540 ;
        RECT  0.180 0.935 0.520 1.275 ;
    END
END OAI2BB1XL

MACRO OAI2BB1X4
    CLASS CORE ;
    FOREIGN OAI2BB1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB1XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.940 0.715 6.120 1.055 ;
        RECT  5.800 0.715 5.940 2.610 ;
        RECT  5.725 0.715 5.800 3.780 ;
        RECT  5.710 0.770 5.725 3.780 ;
        RECT  4.840 0.770 5.710 1.000 ;
        RECT  5.420 2.380 5.710 3.780 ;
        RECT  4.175 2.945 5.420 3.175 ;
        RECT  4.800 0.715 4.840 1.000 ;
        RECT  4.460 0.715 4.800 1.055 ;
        RECT  3.725 2.890 4.175 3.230 ;
        RECT  2.855 2.945 3.725 3.175 ;
        RECT  2.785 2.945 2.855 3.230 ;
        RECT  2.445 2.890 2.785 3.230 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.265 3.020 2.660 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.020 0.520 2.660 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 2.265 1.840 2.660 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 -0.400 6.600 0.400 ;
        RECT  2.740 -0.400 3.080 0.955 ;
        RECT  1.800 -0.400 2.740 0.400 ;
        RECT  1.460 -0.400 1.800 0.955 ;
        RECT  0.000 -0.400 1.460 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.705 4.640 6.600 5.440 ;
        RECT  4.365 3.620 4.705 5.440 ;
        RECT  3.425 4.640 4.365 5.440 ;
        RECT  3.085 3.620 3.425 5.440 ;
        RECT  2.080 4.640 3.085 5.440 ;
        RECT  1.740 3.900 2.080 5.440 ;
        RECT  0.520 4.640 1.740 5.440 ;
        RECT  0.180 3.075 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.140 1.340 5.480 1.780 ;
        RECT  3.905 2.205 5.185 2.545 ;
        RECT  3.840 1.340 5.140 1.570 ;
        RECT  3.565 2.205 3.905 2.435 ;
        RECT  3.500 1.175 3.840 1.570 ;
        RECT  3.335 1.805 3.565 2.435 ;
        RECT  2.385 1.340 3.500 1.570 ;
        RECT  0.980 1.805 3.335 2.035 ;
        RECT  2.155 1.340 2.385 1.575 ;
        RECT  2.100 1.345 2.155 1.575 ;
        RECT  0.980 3.075 1.280 4.355 ;
        RECT  0.940 1.215 0.980 4.355 ;
        RECT  0.750 1.215 0.940 3.310 ;
        RECT  0.520 1.215 0.750 1.445 ;
        RECT  0.180 0.635 0.520 1.445 ;
    END
END OAI2BB1X4

MACRO OAI2BB1X2
    CLASS CORE ;
    FOREIGN OAI2BB1X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB1XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 1.225 3.745 2.635 ;
        RECT  3.515 1.225 3.670 3.070 ;
        RECT  3.160 1.225 3.515 1.455 ;
        RECT  3.440 2.405 3.515 3.070 ;
        RECT  3.260 2.840 3.440 3.070 ;
        RECT  2.920 2.840 3.260 3.180 ;
        RECT  2.820 1.115 3.160 1.455 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.590 2.500 2.130 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.215 1.680 0.585 2.240 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.380 2.020 2.660 ;
        RECT  1.275 2.275 1.505 2.660 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 -0.400 4.620 0.400 ;
        RECT  4.100 -0.400 4.440 1.275 ;
        RECT  1.840 -0.400 4.100 0.400 ;
        RECT  1.500 -0.400 1.840 1.275 ;
        RECT  0.000 -0.400 1.500 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.940 4.640 4.620 5.440 ;
        RECT  3.600 4.465 3.940 5.440 ;
        RECT  2.620 4.640 3.600 5.440 ;
        RECT  2.280 4.020 2.620 5.440 ;
        RECT  1.060 4.640 2.280 5.440 ;
        RECT  0.720 4.465 1.060 5.440 ;
        RECT  0.000 4.640 0.720 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.960 1.965 3.070 2.305 ;
        RECT  2.730 1.965 2.960 2.610 ;
        RECT  2.685 2.380 2.730 2.610 ;
        RECT  2.455 2.380 2.685 3.455 ;
        RECT  1.860 3.225 2.455 3.455 ;
        RECT  1.520 3.225 1.860 3.565 ;
        RECT  1.045 3.225 1.520 3.455 ;
        RECT  0.815 1.175 1.045 3.455 ;
        RECT  0.520 1.175 0.815 1.405 ;
        RECT  0.180 1.065 0.520 1.405 ;
    END
END OAI2BB1X2

MACRO OAI2BB1X1
    CLASS CORE ;
    FOREIGN OAI2BB1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB1XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.440 3.155 3.835 ;
        RECT  2.780 1.440 2.925 1.780 ;
        RECT  2.855 3.525 2.925 3.835 ;
        RECT  2.485 3.605 2.855 3.835 ;
        RECT  2.145 3.605 2.485 3.945 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.210 2.075 2.690 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.570 0.680 2.910 ;
        RECT  0.140 2.570 0.520 3.220 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.625 1.780 1.180 2.235 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.880 -0.400 3.300 0.400 ;
        RECT  1.540 -0.400 1.880 0.575 ;
        RECT  0.000 -0.400 1.540 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.045 4.640 3.300 5.440 ;
        RECT  2.990 4.465 3.045 5.440 ;
        RECT  2.760 4.410 2.990 5.440 ;
        RECT  2.705 4.465 2.760 5.440 ;
        RECT  1.720 4.640 2.705 5.440 ;
        RECT  0.180 4.465 1.720 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.550 2.100 2.695 2.450 ;
        RECT  2.320 0.985 2.550 3.375 ;
        RECT  0.520 0.985 2.320 1.215 ;
        RECT  1.120 3.145 2.320 3.375 ;
        RECT  0.780 3.145 1.120 3.540 ;
        RECT  0.180 0.935 0.520 1.275 ;
    END
END OAI2BB1X1

MACRO OAI22XL
    CLASS CORE ;
    FOREIGN OAI22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.625 3.745 3.755 ;
        RECT  2.910 1.625 3.515 1.855 ;
        RECT  1.840 3.525 3.515 3.755 ;
        RECT  2.760 1.305 2.910 1.855 ;
        RECT  2.680 1.195 2.760 1.855 ;
        RECT  2.420 1.195 2.680 1.535 ;
        RECT  1.500 3.470 1.840 3.810 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.685 0.855 3.220 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.765 1.600 2.130 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.455 3.160 3.220 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.410 2.405 2.425 2.635 ;
        RECT  2.070 1.985 2.410 2.740 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 -0.400 3.960 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 4.640 3.960 5.440 ;
        RECT  2.820 4.465 3.160 5.440 ;
        RECT  0.520 4.640 2.820 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.370 1.055 3.480 1.395 ;
        RECT  3.140 0.735 3.370 1.395 ;
        RECT  2.040 0.735 3.140 0.965 ;
        RECT  1.810 0.735 2.040 1.535 ;
        RECT  1.700 1.195 1.810 1.535 ;
        RECT  0.180 1.250 1.700 1.480 ;
    END
END OAI22XL

MACRO OAI22X4
    CLASS CORE ;
    FOREIGN OAI22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI22XL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.020 1.820 9.100 3.220 ;
        RECT  8.790 0.665 9.020 3.220 ;
        RECT  4.900 0.665 8.790 0.895 ;
        RECT  8.720 1.820 8.790 3.220 ;
        RECT  8.240 2.950 8.720 3.180 ;
        RECT  7.900 2.950 8.240 3.895 ;
        RECT  7.705 2.950 7.900 3.220 ;
        RECT  5.680 2.950 7.705 3.180 ;
        RECT  5.340 2.950 5.680 3.895 ;
        RECT  5.065 2.950 5.340 3.220 ;
        RECT  3.120 2.950 5.065 3.180 ;
        RECT  2.780 2.950 3.120 3.895 ;
        RECT  0.560 2.950 2.780 3.180 ;
        RECT  0.220 2.950 0.560 3.890 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.815 2.255 4.045 2.685 ;
        RECT  2.095 2.455 3.815 2.685 ;
        RECT  1.760 2.310 2.095 2.685 ;
        RECT  1.535 2.310 1.760 2.635 ;
        RECT  1.260 2.310 1.535 2.540 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.810 1.885 3.400 2.225 ;
        RECT  2.540 1.850 2.810 2.225 ;
        RECT  0.445 1.850 2.540 2.080 ;
        RECT  0.215 1.850 0.445 2.635 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.050 1.885 7.160 2.225 ;
        RECT  6.820 1.850 7.050 2.225 ;
        RECT  5.000 1.850 6.820 2.080 ;
        RECT  5.000 2.365 5.065 2.635 ;
        RECT  4.835 1.850 5.000 2.635 ;
        RECT  4.770 1.850 4.835 2.595 ;
        RECT  4.430 2.255 4.770 2.595 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.825 2.255 8.055 2.685 ;
        RECT  7.705 2.380 7.825 2.685 ;
        RECT  6.460 2.455 7.705 2.685 ;
        RECT  6.230 2.310 6.460 2.685 ;
        RECT  6.155 2.310 6.230 2.635 ;
        RECT  5.520 2.310 6.155 2.540 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.800 -0.400 9.240 0.400 ;
        RECT  3.460 -0.400 3.800 0.950 ;
        RECT  2.520 -0.400 3.460 0.400 ;
        RECT  2.180 -0.400 2.520 0.950 ;
        RECT  1.240 -0.400 2.180 0.400 ;
        RECT  0.900 -0.400 1.240 0.950 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.960 4.640 9.240 5.440 ;
        RECT  6.620 3.850 6.960 5.440 ;
        RECT  4.400 4.640 6.620 5.440 ;
        RECT  4.060 3.850 4.400 5.440 ;
        RECT  1.840 4.640 4.060 5.440 ;
        RECT  1.500 3.850 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.220 1.130 8.560 1.470 ;
        RECT  7.690 1.240 8.220 1.470 ;
        RECT  7.460 1.240 7.690 1.620 ;
        RECT  4.520 1.390 7.460 1.620 ;
        RECT  4.180 0.910 4.520 1.620 ;
        RECT  0.965 1.390 4.180 1.620 ;
        RECT  0.735 1.385 0.965 1.620 ;
        RECT  0.520 1.385 0.735 1.615 ;
        RECT  0.290 0.910 0.520 1.615 ;
        RECT  0.180 0.910 0.290 1.250 ;
    END
END OAI22X4

MACRO OAI22X2
    CLASS CORE ;
    FOREIGN OAI22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI22XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.555 1.210 5.785 3.500 ;
        RECT  5.200 1.210 5.555 1.440 ;
        RECT  5.350 3.025 5.555 3.500 ;
        RECT  5.065 3.135 5.350 3.500 ;
        RECT  4.860 1.100 5.200 1.440 ;
        RECT  4.760 3.135 5.065 3.755 ;
        RECT  3.880 1.210 4.860 1.440 ;
        RECT  3.130 3.135 4.760 3.365 ;
        RECT  3.540 1.100 3.880 1.440 ;
        RECT  2.790 3.025 3.130 3.365 ;
        RECT  0.520 3.135 2.790 3.365 ;
        RECT  0.180 3.025 0.520 3.365 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 2.135 2.070 2.475 ;
        RECT  1.105 2.245 1.260 2.475 ;
        RECT  0.875 2.245 1.105 2.635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.685 1.985 2.800 2.325 ;
        RECT  2.460 1.670 2.685 2.325 ;
        RECT  2.455 1.670 2.460 2.270 ;
        RECT  0.520 1.670 2.455 1.900 ;
        RECT  0.180 1.670 0.520 2.325 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.730 4.600 2.325 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.450 5.325 2.790 ;
        RECT  3.745 2.560 4.985 2.790 ;
        RECT  3.520 2.405 3.745 2.790 ;
        RECT  3.130 2.350 3.520 2.790 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 -0.400 5.940 0.400 ;
        RECT  2.060 -0.400 2.400 0.575 ;
        RECT  0.600 -0.400 2.060 0.400 ;
        RECT  0.260 -0.400 0.600 0.575 ;
        RECT  0.000 -0.400 0.260 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 4.640 5.940 5.440 ;
        RECT  4.070 3.765 4.410 5.440 ;
        RECT  1.840 4.640 4.070 5.440 ;
        RECT  1.500 3.765 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.820 1.095 3.160 1.435 ;
        RECT  1.840 1.205 2.820 1.435 ;
        RECT  1.500 1.095 1.840 1.435 ;
        RECT  0.520 1.205 1.500 1.435 ;
        RECT  0.180 1.095 0.520 1.435 ;
    END
END OAI22X2

MACRO OAI22X1
    CLASS CORE ;
    FOREIGN OAI22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI22XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.505 3.745 3.755 ;
        RECT  3.440 1.505 3.515 1.845 ;
        RECT  1.840 3.525 3.515 3.755 ;
        RECT  2.760 1.505 3.440 1.735 ;
        RECT  2.530 1.315 2.760 1.735 ;
        RECT  2.420 1.315 2.530 1.655 ;
        RECT  1.500 3.470 1.840 3.810 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.840 2.750 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.820 1.600 2.185 ;
        RECT  0.800 1.820 1.260 2.145 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.455 3.160 3.220 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.070 1.985 2.500 2.660 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 -0.400 3.960 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 4.640 3.960 5.440 ;
        RECT  2.820 4.465 3.160 5.440 ;
        RECT  0.520 4.640 2.820 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.370 0.935 3.480 1.275 ;
        RECT  3.140 0.855 3.370 1.275 ;
        RECT  2.040 0.855 3.140 1.085 ;
        RECT  1.810 0.855 2.040 1.590 ;
        RECT  1.700 1.250 1.810 1.590 ;
        RECT  0.520 1.305 1.700 1.535 ;
        RECT  0.180 1.250 0.520 1.590 ;
    END
END OAI22X1

MACRO OAI222XL
    CLASS CORE ;
    FOREIGN OAI222XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.760 5.065 3.755 ;
        RECT  4.480 1.760 4.835 1.990 ;
        RECT  4.330 3.525 4.835 3.755 ;
        RECT  4.340 1.515 4.480 1.990 ;
        RECT  4.110 1.180 4.340 1.990 ;
        RECT  3.990 3.480 4.330 3.820 ;
        RECT  4.000 1.180 4.110 1.520 ;
        RECT  3.745 3.500 3.990 3.780 ;
        RECT  1.640 3.535 3.745 3.765 ;
        RECT  1.300 3.480 1.640 3.820 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.245 2.130 3.820 2.660 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.095 2.585 4.580 3.220 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.520 3.005 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.735 1.270 2.345 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.425 2.550 3.225 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 2.685 1.840 3.220 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 5.280 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.985 4.640 5.280 5.440 ;
        RECT  2.645 4.465 2.985 5.440 ;
        RECT  0.520 4.640 2.645 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.950 1.180 5.060 1.520 ;
        RECT  4.720 0.650 4.950 1.520 ;
        RECT  3.620 0.650 4.720 0.880 ;
        RECT  3.390 0.650 3.620 1.520 ;
        RECT  3.280 1.180 3.390 1.520 ;
        RECT  2.560 1.060 2.900 1.520 ;
        RECT  1.080 1.060 2.560 1.290 ;
        RECT  0.740 1.060 1.080 1.400 ;
    END
END OAI222XL

MACRO OAI222X4
    CLASS CORE ;
    FOREIGN OAI222X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI222XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.970 1.820 7.120 3.220 ;
        RECT  6.920 1.500 6.970 3.220 ;
        RECT  6.905 0.920 6.920 3.220 ;
        RECT  6.740 0.920 6.905 4.170 ;
        RECT  6.580 0.920 6.740 1.730 ;
        RECT  6.565 2.890 6.740 4.170 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.145 3.820 2.780 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 2.380 4.480 3.105 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.520 2.510 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.655 2.770 1.270 3.395 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 2.765 3.160 3.245 ;
        RECT  2.455 2.765 2.460 3.105 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 1.820 2.185 2.465 ;
        RECT  1.780 1.820 2.120 2.470 ;
        RECT  1.460 1.820 1.780 2.465 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.640 -0.400 7.920 0.400 ;
        RECT  7.300 -0.400 7.640 1.425 ;
        RECT  6.200 -0.400 7.300 0.400 ;
        RECT  5.860 -0.400 6.200 0.950 ;
        RECT  1.640 -0.400 5.860 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.625 4.640 7.920 5.440 ;
        RECT  7.285 3.620 7.625 5.440 ;
        RECT  6.145 4.640 7.285 5.440 ;
        RECT  5.805 4.465 6.145 5.440 ;
        RECT  4.825 4.640 5.805 5.440 ;
        RECT  4.485 4.465 4.825 5.440 ;
        RECT  2.965 4.640 4.485 5.440 ;
        RECT  2.625 4.465 2.965 5.440 ;
        RECT  0.520 4.640 2.625 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.160 2.250 6.500 2.590 ;
        RECT  5.810 2.305 6.160 2.590 ;
        RECT  5.580 1.260 5.810 3.930 ;
        RECT  5.480 1.260 5.580 1.490 ;
        RECT  5.245 3.590 5.580 3.930 ;
        RECT  5.140 0.680 5.480 1.490 ;
        RECT  4.945 2.470 5.345 2.810 ;
        RECT  4.715 1.920 4.945 3.870 ;
        RECT  4.280 1.920 4.715 2.150 ;
        RECT  4.325 3.640 4.715 3.870 ;
        RECT  3.985 3.640 4.325 3.980 ;
        RECT  4.050 1.420 4.280 2.150 ;
        RECT  3.880 1.420 4.050 1.760 ;
        RECT  1.640 3.640 3.985 3.870 ;
        RECT  2.560 1.250 2.900 1.760 ;
        RECT  1.080 1.250 2.560 1.480 ;
        RECT  1.300 3.640 1.640 3.980 ;
        RECT  0.740 1.140 1.080 1.480 ;
    END
END OAI222X4

MACRO OAI222X2
    CLASS CORE ;
    FOREIGN OAI222X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI222XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.660 1.390 8.890 3.730 ;
        RECT  7.085 1.390 8.660 1.620 ;
        RECT  8.365 3.500 8.660 3.730 ;
        RECT  8.135 3.500 8.365 3.755 ;
        RECT  7.480 3.525 8.135 3.755 ;
        RECT  7.040 3.525 7.480 3.865 ;
        RECT  4.840 3.525 7.040 3.755 ;
        RECT  4.395 3.525 4.840 3.865 ;
        RECT  2.240 3.525 4.395 3.755 ;
        RECT  1.900 3.525 2.240 3.865 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.320 2.835 8.430 3.065 ;
        RECT  8.090 2.835 8.320 3.120 ;
        RECT  6.600 2.890 8.090 3.120 ;
        RECT  6.370 2.405 6.600 3.120 ;
        RECT  6.155 2.405 6.370 2.635 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.400 2.090 7.780 2.660 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.320 3.150 2.550 ;
        RECT  0.920 2.320 1.105 2.635 ;
        RECT  0.580 2.295 0.920 2.635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.780 2.480 3.120 ;
        RECT  2.195 2.780 2.425 3.195 ;
        RECT  1.660 2.780 2.195 3.120 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.415 2.360 5.845 2.590 ;
        RECT  5.185 2.320 5.415 2.590 ;
        RECT  4.000 2.320 5.185 2.550 ;
        RECT  3.770 2.320 4.000 2.690 ;
        RECT  3.660 2.350 3.770 2.690 ;
        RECT  3.515 2.405 3.660 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.940 2.940 5.105 3.220 ;
        RECT  4.600 2.780 4.940 3.220 ;
        RECT  4.300 2.940 4.600 3.220 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 -0.400 9.900 0.400 ;
        RECT  2.900 -0.400 3.240 0.950 ;
        RECT  1.800 -0.400 2.900 0.400 ;
        RECT  1.460 -0.400 1.800 0.950 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.680 4.640 9.900 5.440 ;
        RECT  8.340 4.070 8.680 5.440 ;
        RECT  6.080 4.640 8.340 5.440 ;
        RECT  5.740 4.070 6.080 5.440 ;
        RECT  3.520 4.640 5.740 5.440 ;
        RECT  3.180 4.070 3.520 5.440 ;
        RECT  0.960 4.640 3.180 5.440 ;
        RECT  0.620 4.070 0.960 5.440 ;
        RECT  0.000 4.640 0.620 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.650 0.810 9.470 1.040 ;
        RECT  6.420 0.665 6.650 1.375 ;
        RECT  3.600 0.665 6.420 0.895 ;
        RECT  4.580 1.270 5.985 1.500 ;
        RECT  4.240 1.270 4.580 1.675 ;
        RECT  2.520 1.270 4.240 1.500 ;
        RECT  2.410 0.890 2.520 1.500 ;
        RECT  2.180 0.890 2.410 1.565 ;
        RECT  1.160 1.335 2.180 1.565 ;
        RECT  0.820 1.335 1.160 1.675 ;
    END
END OAI222X2

MACRO OAI222X1
    CLASS CORE ;
    FOREIGN OAI222X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI222XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.600 3.480 5.780 3.820 ;
        RECT  5.370 1.515 5.600 3.820 ;
        RECT  4.880 1.515 5.370 1.745 ;
        RECT  2.170 3.480 5.370 3.820 ;
        RECT  4.540 1.405 4.880 1.745 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.985 4.480 2.660 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.760 2.455 5.140 3.220 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.840 2.750 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.695 1.880 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.425 3.550 2.970 ;
        RECT  3.210 2.425 3.440 3.170 ;
        RECT  3.085 2.940 3.210 3.170 ;
        RECT  2.855 2.940 3.085 3.195 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 2.380 2.880 2.660 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 -0.400 5.940 0.400 ;
        RECT  1.700 -0.400 2.040 0.575 ;
        RECT  0.520 -0.400 1.700 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.830 4.640 5.940 5.440 ;
        RECT  3.490 4.465 3.830 5.440 ;
        RECT  1.190 4.640 3.490 5.440 ;
        RECT  1.135 4.465 1.190 5.440 ;
        RECT  0.905 4.410 1.135 5.440 ;
        RECT  0.850 4.465 0.905 5.440 ;
        RECT  0.000 4.640 0.850 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.260 0.920 5.600 1.260 ;
        RECT  4.160 0.940 5.260 1.170 ;
        RECT  4.050 0.940 4.160 1.280 ;
        RECT  3.820 0.940 4.050 1.715 ;
        RECT  2.380 1.485 3.820 1.715 ;
        RECT  1.280 1.005 3.440 1.235 ;
        RECT  0.940 0.895 1.280 1.235 ;
    END
END OAI222X1

MACRO OAI221XL
    CLASS CORE ;
    FOREIGN OAI221XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.085 4.405 3.865 ;
        RECT  3.890 1.085 4.175 1.425 ;
        RECT  3.520 3.635 4.175 3.865 ;
        RECT  3.180 3.635 3.520 3.975 ;
        RECT  1.640 3.635 3.180 3.865 ;
        RECT  1.300 3.635 1.640 3.975 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.190 3.820 2.745 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.690 0.520 3.450 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.665 1.820 1.275 2.310 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 2.940 3.085 3.195 ;
        RECT  2.550 2.940 2.855 3.170 ;
        RECT  2.210 2.685 2.550 3.170 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.835 2.695 1.845 3.270 ;
        RECT  1.495 2.690 1.835 3.270 ;
        RECT  1.195 2.695 1.495 3.270 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 4.620 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 4.640 4.620 5.440 ;
        RECT  2.420 4.465 2.760 5.440 ;
        RECT  0.520 4.640 2.420 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.795 1.425 2.905 1.765 ;
        RECT  2.565 1.060 2.795 1.765 ;
        RECT  1.080 1.060 2.565 1.290 ;
        RECT  0.740 1.060 1.080 1.400 ;
    END
END OAI221XL

MACRO OAI221X4
    CLASS CORE ;
    FOREIGN OAI221X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI221XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.820 6.460 3.220 ;
        RECT  6.200 1.220 6.315 3.220 ;
        RECT  6.105 0.645 6.200 3.220 ;
        RECT  6.085 0.645 6.105 4.095 ;
        RECT  5.860 0.645 6.085 1.455 ;
        RECT  6.080 1.820 6.085 4.095 ;
        RECT  5.765 2.815 6.080 4.095 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 2.350 3.820 2.925 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.745 0.600 3.320 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.710 1.470 2.170 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 2.405 3.085 2.660 ;
        RECT  2.555 2.430 2.855 2.660 ;
        RECT  2.325 2.430 2.555 3.085 ;
        RECT  2.215 2.745 2.325 3.085 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.735 1.880 3.315 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.920 -0.400 7.260 0.400 ;
        RECT  6.580 -0.400 6.920 1.420 ;
        RECT  5.480 -0.400 6.580 0.400 ;
        RECT  5.140 -0.400 5.480 1.425 ;
        RECT  1.640 -0.400 5.140 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.825 4.640 7.260 5.440 ;
        RECT  6.485 3.615 6.825 5.440 ;
        RECT  5.345 4.640 6.485 5.440 ;
        RECT  5.005 4.465 5.345 5.440 ;
        RECT  4.225 4.640 5.005 5.440 ;
        RECT  3.885 4.465 4.225 5.440 ;
        RECT  2.760 4.640 3.885 5.440 ;
        RECT  2.420 4.465 2.760 5.440 ;
        RECT  0.520 4.640 2.420 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.355 1.920 5.695 2.260 ;
        RECT  5.005 1.975 5.355 2.260 ;
        RECT  4.785 1.690 5.005 3.920 ;
        RECT  4.775 1.690 4.785 3.975 ;
        RECT  4.760 1.690 4.775 1.920 ;
        RECT  4.445 3.635 4.775 3.975 ;
        RECT  4.530 0.905 4.760 1.920 ;
        RECT  4.280 2.285 4.545 2.625 ;
        RECT  4.420 0.905 4.530 1.245 ;
        RECT  4.050 1.615 4.280 3.400 ;
        RECT  3.880 1.615 4.050 1.955 ;
        RECT  3.525 3.170 4.050 3.400 ;
        RECT  3.295 3.170 3.525 3.965 ;
        RECT  1.300 3.625 3.295 3.965 ;
        RECT  2.560 1.250 2.900 1.760 ;
        RECT  1.080 1.250 2.560 1.480 ;
        RECT  0.740 1.140 1.080 1.480 ;
    END
END OAI221X4

MACRO OAI221X2
    CLASS CORE ;
    FOREIGN OAI221X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI221XL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.450 7.580 3.485 ;
        RECT  7.350 1.335 7.370 3.485 ;
        RECT  7.140 1.335 7.350 1.850 ;
        RECT  6.460 3.255 7.350 3.485 ;
        RECT  6.400 3.255 6.460 3.525 ;
        RECT  6.170 3.255 6.400 3.795 ;
        RECT  6.060 3.455 6.170 3.795 ;
        RECT  4.360 3.525 6.060 3.755 ;
        RECT  4.020 3.525 4.360 3.865 ;
        RECT  3.740 3.525 4.020 3.780 ;
        RECT  1.800 3.525 3.740 3.755 ;
        RECT  1.460 3.525 1.800 3.865 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.145 2.380 7.100 2.660 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 2.320 2.760 2.550 ;
        RECT  0.420 2.295 0.760 2.635 ;
        RECT  0.215 2.405 0.420 2.635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 2.780 2.040 3.120 ;
        RECT  1.535 2.780 1.765 3.195 ;
        RECT  1.220 2.780 1.535 3.120 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.920 2.360 5.640 2.590 ;
        RECT  4.690 2.320 4.920 2.590 ;
        RECT  3.745 2.320 4.690 2.550 ;
        RECT  3.560 2.320 3.745 2.635 ;
        RECT  3.515 2.320 3.560 2.690 ;
        RECT  3.220 2.350 3.515 2.690 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.460 2.940 4.625 3.220 ;
        RECT  4.120 2.780 4.460 3.220 ;
        RECT  3.820 2.940 4.120 3.220 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 -0.400 8.580 0.400 ;
        RECT  2.900 -0.400 3.240 0.950 ;
        RECT  1.800 -0.400 2.900 0.400 ;
        RECT  1.460 -0.400 1.800 0.950 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.120 4.640 8.580 5.440 ;
        RECT  6.780 3.715 7.120 5.440 ;
        RECT  5.640 4.640 6.780 5.440 ;
        RECT  5.300 4.070 5.640 5.440 ;
        RECT  3.080 4.640 5.300 5.440 ;
        RECT  2.740 4.070 3.080 5.440 ;
        RECT  0.520 4.640 2.740 5.440 ;
        RECT  0.180 3.840 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.650 0.810 8.065 1.040 ;
        RECT  6.420 0.665 6.650 1.375 ;
        RECT  3.600 0.665 6.420 0.895 ;
        RECT  4.580 1.270 5.985 1.500 ;
        RECT  4.240 1.270 4.580 1.675 ;
        RECT  2.520 1.270 4.240 1.500 ;
        RECT  2.410 0.910 2.520 1.500 ;
        RECT  2.180 0.910 2.410 1.565 ;
        RECT  1.160 1.335 2.180 1.565 ;
        RECT  0.820 1.335 1.160 1.675 ;
    END
END OAI221X2

MACRO OAI221X1
    CLASS CORE ;
    FOREIGN OAI221X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI221XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.940 3.480 5.120 3.820 ;
        RECT  4.710 1.185 4.940 3.820 ;
        RECT  4.540 1.185 4.710 1.525 ;
        RECT  1.500 3.480 4.710 3.820 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.835 2.240 4.480 2.690 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.840 2.750 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.675 1.555 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.540 2.380 3.160 2.820 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.415 2.350 2.190 2.825 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 -0.400 5.280 0.400 ;
        RECT  1.700 -0.400 2.040 0.575 ;
        RECT  0.520 -0.400 1.700 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 4.640 5.280 5.440 ;
        RECT  3.105 4.465 3.160 5.440 ;
        RECT  2.875 4.410 3.105 5.440 ;
        RECT  2.820 4.465 2.875 5.440 ;
        RECT  0.520 4.640 2.820 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.820 1.415 4.160 1.755 ;
        RECT  2.720 1.525 3.820 1.755 ;
        RECT  3.100 0.950 3.440 1.290 ;
        RECT  1.280 0.950 3.100 1.180 ;
        RECT  2.380 1.450 2.720 1.790 ;
        RECT  0.940 0.950 1.280 1.290 ;
    END
END OAI221X1

MACRO OAI21XL
    CLASS CORE ;
    FOREIGN OAI21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.845 2.450 3.845 ;
        RECT  2.220 0.675 2.425 3.845 ;
        RECT  2.195 0.675 2.220 2.075 ;
        RECT  1.800 3.615 2.220 3.845 ;
        RECT  2.060 0.675 2.195 0.905 ;
        RECT  1.460 3.560 1.800 3.900 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.690 1.990 3.220 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.180 1.820 0.520 2.595 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.010 1.465 2.400 ;
        RECT  0.875 1.845 1.105 2.400 ;
        RECT  0.800 2.010 0.875 2.400 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 -0.400 2.640 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 4.640 2.640 5.440 ;
        RECT  2.020 4.465 2.360 5.440 ;
        RECT  0.520 4.640 2.020 5.440 ;
        RECT  0.180 3.760 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.730 1.395 1.840 1.735 ;
        RECT  1.500 1.245 1.730 1.735 ;
        RECT  0.520 1.245 1.500 1.475 ;
        RECT  0.180 1.245 0.520 1.585 ;
    END
END OAI21XL

MACRO OAI21X4
    CLASS CORE ;
    FOREIGN OAI21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI21XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.460 1.315 6.565 1.850 ;
        RECT  6.225 1.315 6.460 3.220 ;
        RECT  6.080 1.390 6.225 3.220 ;
        RECT  4.825 1.390 6.080 1.620 ;
        RECT  5.720 2.975 6.080 3.205 ;
        RECT  5.380 2.920 5.720 3.260 ;
        RECT  4.440 2.975 5.380 3.205 ;
        RECT  4.330 2.920 4.440 3.260 ;
        RECT  4.100 2.920 4.330 3.635 ;
        RECT  1.800 3.405 4.100 3.635 ;
        RECT  1.460 3.350 1.800 3.690 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 2.350 5.400 2.690 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.860 2.310 3.400 2.540 ;
        RECT  2.730 2.310 2.860 2.660 ;
        RECT  2.500 2.310 2.730 3.120 ;
        RECT  0.760 2.890 2.500 3.120 ;
        RECT  0.530 2.240 0.760 3.120 ;
        RECT  0.475 2.240 0.530 2.660 ;
        RECT  0.420 2.240 0.475 2.635 ;
        RECT  0.215 2.405 0.420 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.960 2.120 4.070 2.460 ;
        RECT  3.730 1.850 3.960 2.460 ;
        RECT  2.120 1.850 3.730 2.080 ;
        RECT  1.890 1.850 2.120 2.580 ;
        RECT  1.785 2.240 1.890 2.580 ;
        RECT  1.535 2.240 1.785 2.635 ;
        RECT  1.220 2.240 1.535 2.580 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.800 -0.400 7.260 0.400 ;
        RECT  3.460 -0.400 3.800 0.950 ;
        RECT  2.520 -0.400 3.460 0.400 ;
        RECT  2.180 -0.400 2.520 0.950 ;
        RECT  1.240 -0.400 2.180 0.400 ;
        RECT  0.900 -0.400 1.240 0.950 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.365 4.640 7.260 5.440 ;
        RECT  6.025 3.645 6.365 5.440 ;
        RECT  5.080 4.640 6.025 5.440 ;
        RECT  4.740 3.645 5.080 5.440 ;
        RECT  3.120 4.640 4.740 5.440 ;
        RECT  2.780 3.915 3.120 5.440 ;
        RECT  0.520 4.640 2.780 5.440 ;
        RECT  0.180 3.495 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.465 0.630 5.805 0.970 ;
        RECT  4.525 0.685 5.465 0.915 ;
        RECT  4.415 0.630 4.525 0.970 ;
        RECT  4.185 0.630 4.415 1.620 ;
        RECT  0.520 1.390 4.185 1.620 ;
        RECT  0.290 0.950 0.520 1.620 ;
        RECT  0.180 0.950 0.290 1.290 ;
    END
END OAI21X4

MACRO OAI21X2
    CLASS CORE ;
    FOREIGN OAI21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI21XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.840 1.305 5.065 3.865 ;
        RECT  4.835 1.305 4.840 3.975 ;
        RECT  4.200 1.305 4.835 1.535 ;
        RECT  4.340 3.635 4.835 3.975 ;
        RECT  3.160 3.635 4.340 3.865 ;
        RECT  3.970 1.105 4.200 1.535 ;
        RECT  3.860 1.105 3.970 1.445 ;
        RECT  2.820 3.635 3.160 3.975 ;
        RECT  0.520 3.635 2.820 3.865 ;
        RECT  0.180 3.635 0.520 3.975 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 2.315 4.445 2.655 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 2.580 2.120 2.920 ;
        RECT  1.785 2.580 1.840 2.970 ;
        RECT  1.535 2.580 1.785 3.195 ;
        RECT  1.220 2.580 1.535 2.970 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 2.540 2.790 2.880 ;
        RECT  2.450 1.930 2.680 2.880 ;
        RECT  0.875 1.930 2.450 2.160 ;
        RECT  0.450 1.820 0.875 2.160 ;
        RECT  0.445 1.845 0.450 2.160 ;
        RECT  0.215 1.845 0.445 2.075 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 -0.400 5.280 0.400 ;
        RECT  2.420 -0.400 2.760 1.240 ;
        RECT  1.280 -0.400 2.420 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.920 4.640 5.280 5.440 ;
        RECT  3.580 4.465 3.920 5.440 ;
        RECT  1.840 4.640 3.580 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.810 0.735 4.920 1.075 ;
        RECT  4.580 0.645 4.810 1.075 ;
        RECT  3.480 0.645 4.580 0.875 ;
        RECT  3.370 0.645 3.480 1.190 ;
        RECT  3.250 0.645 3.370 1.700 ;
        RECT  3.140 0.850 3.250 1.700 ;
        RECT  2.040 1.470 3.140 1.700 ;
        RECT  1.985 0.935 2.040 1.700 ;
        RECT  1.810 0.930 1.985 1.700 ;
        RECT  1.700 0.930 1.810 1.275 ;
        RECT  0.520 0.930 1.700 1.160 ;
        RECT  0.180 0.820 0.520 1.160 ;
    END
END OAI21X2

MACRO OAI21X1
    CLASS CORE ;
    FOREIGN OAI21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI21XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.860 1.235 3.085 3.845 ;
        RECT  2.855 1.125 2.860 3.845 ;
        RECT  2.420 1.125 2.855 1.465 ;
        RECT  1.880 3.615 2.855 3.845 ;
        RECT  1.540 3.560 1.880 3.900 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.030 2.350 2.500 2.955 ;
        RECT  2.020 2.350 2.030 2.690 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 1.820 0.880 2.100 ;
        RECT  0.260 1.790 0.600 2.130 ;
        RECT  0.140 1.820 0.260 2.100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.560 2.660 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 -0.400 3.300 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.640 4.640 3.300 5.440 ;
        RECT  2.300 4.465 2.640 5.440 ;
        RECT  0.520 4.640 2.300 5.440 ;
        RECT  0.180 3.740 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.985 0.935 2.040 1.275 ;
        RECT  1.700 0.915 1.985 1.275 ;
        RECT  0.520 0.915 1.700 1.145 ;
        RECT  0.180 0.860 0.520 1.200 ;
    END
END OAI21X1

MACRO OAI211XL
    CLASS CORE ;
    FOREIGN OAI211XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 1.250 3.745 3.790 ;
        RECT  3.515 1.140 3.520 3.900 ;
        RECT  3.020 1.140 3.515 1.480 ;
        RECT  3.060 3.560 3.515 3.900 ;
        RECT  1.880 3.560 3.060 3.790 ;
        RECT  1.540 3.560 1.880 3.900 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.030 2.350 2.500 2.955 ;
        RECT  2.020 2.350 2.030 2.690 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.820 3.160 2.530 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 1.820 0.880 2.100 ;
        RECT  0.260 1.790 0.600 2.130 ;
        RECT  0.140 1.820 0.260 2.100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.560 2.660 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 -0.400 3.960 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.640 4.640 3.960 5.440 ;
        RECT  2.300 4.465 2.640 5.440 ;
        RECT  0.520 4.640 2.300 5.440 ;
        RECT  0.180 3.560 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.700 0.860 2.040 1.200 ;
        RECT  0.520 0.915 1.700 1.145 ;
        RECT  0.180 0.860 0.520 1.200 ;
    END
END OAI211XL

MACRO OAI211X4
    CLASS CORE ;
    FOREIGN OAI211X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI211XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 1.260 5.800 2.660 ;
        RECT  5.420 1.260 5.760 3.180 ;
        RECT  4.780 1.335 5.420 1.675 ;
        RECT  4.460 2.840 5.420 3.180 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.370 1.790 2.080 2.130 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 2.255 3.160 2.780 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 2.390 1.360 2.730 ;
        RECT  1.020 2.390 1.250 3.195 ;
        RECT  0.875 2.965 1.020 3.195 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.145 0.690 2.665 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 -0.400 5.940 0.400 ;
        RECT  5.420 -0.400 5.760 0.950 ;
        RECT  4.480 -0.400 5.420 0.400 ;
        RECT  4.140 -0.400 4.480 0.950 ;
        RECT  1.180 -0.400 4.140 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.440 4.640 5.940 5.440 ;
        RECT  5.100 4.020 5.440 5.440 ;
        RECT  4.160 4.640 5.100 5.440 ;
        RECT  3.820 4.020 4.160 5.440 ;
        RECT  2.600 4.640 3.820 5.440 ;
        RECT  1.500 4.465 2.600 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.230 1.940 4.980 2.280 ;
        RECT  4.000 1.180 4.230 3.790 ;
        RECT  3.720 1.180 4.000 1.410 ;
        RECT  3.400 3.560 4.000 3.790 ;
        RECT  3.660 2.030 3.770 2.370 ;
        RECT  3.490 0.630 3.720 1.410 ;
        RECT  3.430 1.655 3.660 3.330 ;
        RECT  3.380 0.630 3.490 0.970 ;
        RECT  3.160 1.655 3.430 1.885 ;
        RECT  2.400 3.100 3.430 3.330 ;
        RECT  3.060 3.560 3.400 3.900 ;
        RECT  2.930 1.330 3.160 1.885 ;
        RECT  2.820 1.330 2.930 1.670 ;
        RECT  2.290 3.100 2.400 3.440 ;
        RECT  2.060 3.100 2.290 3.920 ;
        RECT  0.520 3.690 2.060 3.920 ;
        RECT  1.500 1.130 1.840 1.470 ;
        RECT  0.520 1.165 1.500 1.395 ;
        RECT  0.180 1.080 0.520 1.420 ;
        RECT  0.180 3.690 0.520 4.030 ;
    END
END OAI211X4

MACRO OAI211X2
    CLASS CORE ;
    FOREIGN OAI211X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI211XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 1.300 6.210 3.170 ;
        RECT  4.835 1.300 5.980 1.530 ;
        RECT  5.725 2.940 5.980 3.170 ;
        RECT  5.650 2.940 5.725 3.195 ;
        RECT  5.495 2.940 5.650 3.865 ;
        RECT  5.420 2.965 5.495 3.865 ;
        RECT  4.840 3.635 5.420 3.865 ;
        RECT  4.340 3.635 4.840 3.975 ;
        RECT  4.760 1.285 4.835 1.530 ;
        RECT  4.420 1.190 4.760 1.530 ;
        RECT  3.160 3.635 4.340 3.865 ;
        RECT  2.820 3.635 3.160 4.000 ;
        RECT  0.520 3.635 2.820 3.865 ;
        RECT  0.180 3.635 0.520 3.975 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.640 1.760 5.750 2.100 ;
        RECT  5.410 1.760 5.640 2.635 ;
        RECT  3.715 2.405 5.410 2.635 ;
        RECT  3.485 1.930 3.715 2.635 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.000 1.845 5.065 2.075 ;
        RECT  4.180 1.790 5.000 2.130 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 2.580 2.120 2.920 ;
        RECT  1.785 2.580 1.840 2.970 ;
        RECT  1.535 2.580 1.785 3.195 ;
        RECT  1.220 2.580 1.535 2.970 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 2.540 2.790 2.880 ;
        RECT  2.450 1.930 2.680 2.880 ;
        RECT  0.875 1.930 2.450 2.160 ;
        RECT  0.790 1.820 0.875 2.160 ;
        RECT  0.450 1.790 0.790 2.160 ;
        RECT  0.445 1.845 0.450 2.160 ;
        RECT  0.215 1.845 0.445 2.075 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 -0.400 6.600 0.400 ;
        RECT  2.420 -0.400 2.760 1.240 ;
        RECT  1.280 -0.400 2.420 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.920 4.640 6.600 5.440 ;
        RECT  3.580 4.465 3.920 5.440 ;
        RECT  1.840 4.640 3.580 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.700 0.720 6.040 1.060 ;
        RECT  3.480 0.730 5.700 0.960 ;
        RECT  3.370 0.730 3.480 1.190 ;
        RECT  3.250 0.730 3.370 1.700 ;
        RECT  3.140 0.850 3.250 1.700 ;
        RECT  2.040 1.470 3.140 1.700 ;
        RECT  1.985 0.935 2.040 1.700 ;
        RECT  1.810 0.930 1.985 1.700 ;
        RECT  1.700 0.930 1.810 1.275 ;
        RECT  0.520 0.930 1.700 1.160 ;
        RECT  0.180 0.820 0.520 1.160 ;
    END
END OAI211X2

MACRO OAI211X1
    CLASS CORE ;
    FOREIGN OAI211X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI211XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 1.250 3.745 3.790 ;
        RECT  3.515 1.140 3.520 3.900 ;
        RECT  3.020 1.140 3.515 1.480 ;
        RECT  3.060 3.560 3.515 3.900 ;
        RECT  1.880 3.560 3.060 3.790 ;
        RECT  1.540 3.560 1.880 3.900 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.030 2.350 2.500 2.955 ;
        RECT  2.020 2.350 2.030 2.690 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.820 3.160 2.530 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 1.820 0.880 2.100 ;
        RECT  0.260 1.790 0.600 2.130 ;
        RECT  0.140 1.820 0.260 2.100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.560 2.660 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 -0.400 3.960 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.640 4.640 3.960 5.440 ;
        RECT  2.300 4.465 2.640 5.440 ;
        RECT  0.520 4.640 2.300 5.440 ;
        RECT  0.180 3.740 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.700 0.860 2.040 1.200 ;
        RECT  0.520 0.915 1.700 1.145 ;
        RECT  0.180 0.860 0.520 1.200 ;
    END
END OAI211X1

MACRO NOR4BBXL
    CLASS CORE ;
    FOREIGN NOR4BBXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.930 0.805 5.160 3.755 ;
        RECT  3.355 0.805 4.930 1.035 ;
        RECT  3.825 3.525 4.930 3.755 ;
        RECT  3.485 3.525 3.825 3.865 ;
        RECT  3.350 0.805 3.355 1.400 ;
        RECT  3.125 0.805 3.350 1.455 ;
        RECT  1.575 1.115 3.125 1.455 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.520 2.405 1.765 2.635 ;
        RECT  1.290 1.690 1.520 2.635 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 2.405 2.425 2.635 ;
        RECT  2.110 1.730 2.340 2.635 ;
        RECT  1.905 1.730 2.110 2.070 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 2.275 4.205 2.615 ;
        RECT  3.855 2.275 4.085 3.195 ;
        RECT  3.515 2.940 3.855 3.195 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.175 1.840 0.515 2.500 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 -0.400 5.280 0.400 ;
        RECT  3.770 -0.400 4.110 0.575 ;
        RECT  2.770 -0.400 3.770 0.400 ;
        RECT  2.430 -0.400 2.770 0.575 ;
        RECT  1.155 -0.400 2.430 0.400 ;
        RECT  0.815 -0.400 1.155 0.575 ;
        RECT  0.000 -0.400 0.815 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.655 4.640 5.280 5.440 ;
        RECT  4.315 4.015 4.655 5.440 ;
        RECT  1.270 4.640 4.315 5.440 ;
        RECT  0.930 4.410 1.270 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.455 1.265 4.685 3.270 ;
        RECT  2.915 1.780 4.455 2.010 ;
        RECT  4.315 2.930 4.455 3.270 ;
        RECT  3.245 2.275 3.585 2.620 ;
        RECT  3.005 2.390 3.245 2.620 ;
        RECT  2.775 2.390 3.005 3.125 ;
        RECT  2.575 1.780 2.915 2.160 ;
        RECT  0.990 2.895 2.775 3.125 ;
        RECT  0.760 1.225 0.990 3.125 ;
        RECT  0.520 1.225 0.760 1.455 ;
        RECT  0.520 2.805 0.760 3.125 ;
        RECT  0.180 1.115 0.520 1.455 ;
        RECT  0.180 2.805 0.520 3.145 ;
    END
END NOR4BBXL

MACRO NOR4BBX4
    CLASS CORE ;
    FOREIGN NOR4BBX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BBXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.990 2.380 13.060 3.780 ;
        RECT  12.760 0.980 12.990 3.780 ;
        RECT  11.960 0.980 12.760 1.210 ;
        RECT  12.680 2.380 12.760 3.780 ;
        RECT  8.885 3.550 12.680 3.780 ;
        RECT  11.730 0.980 11.960 1.415 ;
        RECT  10.780 1.185 11.730 1.415 ;
        RECT  10.440 1.075 10.780 1.415 ;
        RECT  9.340 1.185 10.440 1.415 ;
        RECT  9.000 1.075 9.340 1.415 ;
        RECT  3.400 1.185 9.000 1.415 ;
        RECT  8.545 3.550 8.885 4.235 ;
        RECT  3.825 4.005 8.545 4.235 ;
        RECT  3.485 4.005 3.825 4.345 ;
        RECT  3.060 1.075 3.400 1.415 ;
        RECT  1.960 1.185 3.060 1.415 ;
        RECT  1.620 1.075 1.960 1.415 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.795 2.195 11.080 3.185 ;
        RECT  6.385 2.955 10.795 3.185 ;
        RECT  6.330 2.955 6.385 3.195 ;
        RECT  6.220 2.595 6.330 3.195 ;
        RECT  5.990 2.595 6.220 3.775 ;
        RECT  1.535 3.545 5.990 3.775 ;
        RECT  1.520 3.500 1.535 3.775 ;
        RECT  1.290 2.210 1.520 3.775 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.355 2.195 10.465 2.535 ;
        RECT  10.125 2.195 10.355 2.720 ;
        RECT  7.220 2.490 10.125 2.720 ;
        RECT  6.990 2.110 7.220 2.720 ;
        RECT  6.740 2.110 6.990 2.450 ;
        RECT  5.490 2.110 6.740 2.340 ;
        RECT  5.380 2.110 5.490 2.450 ;
        RECT  5.140 2.110 5.380 3.315 ;
        RECT  4.835 2.965 5.140 3.315 ;
        RECT  2.245 3.085 4.835 3.315 ;
        RECT  2.015 2.335 2.245 3.315 ;
        RECT  1.905 2.335 2.015 2.675 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.380 2.120 11.945 2.645 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.170 1.845 0.510 2.555 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.500 -0.400 13.200 0.400 ;
        RECT  11.160 -0.400 11.500 0.955 ;
        RECT  10.060 -0.400 11.160 0.400 ;
        RECT  9.720 -0.400 10.060 0.955 ;
        RECT  8.620 -0.400 9.720 0.400 ;
        RECT  8.280 -0.400 8.620 0.955 ;
        RECT  4.135 -0.400 8.280 0.400 ;
        RECT  3.795 -0.400 4.135 0.955 ;
        RECT  2.680 -0.400 3.795 0.400 ;
        RECT  2.340 -0.400 2.680 0.950 ;
        RECT  1.240 -0.400 2.340 0.400 ;
        RECT  0.900 -0.400 1.240 0.950 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.530 4.640 13.200 5.440 ;
        RECT  11.190 4.465 11.530 5.440 ;
        RECT  6.355 4.640 11.190 5.440 ;
        RECT  6.015 4.465 6.355 5.440 ;
        RECT  1.295 4.640 6.015 5.440 ;
        RECT  0.955 4.465 1.295 5.440 ;
        RECT  0.000 4.640 0.955 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.435 1.450 12.530 1.880 ;
        RECT  12.205 1.450 12.435 3.230 ;
        RECT  12.190 1.450 12.205 1.875 ;
        RECT  11.950 2.890 12.205 3.230 ;
        RECT  9.795 1.645 12.190 1.875 ;
        RECT  9.565 1.645 9.795 2.260 ;
        RECT  9.455 1.920 9.565 2.260 ;
        RECT  7.970 2.030 9.455 2.260 ;
        RECT  7.860 1.920 7.970 2.260 ;
        RECT  7.630 1.645 7.860 2.260 ;
        RECT  4.740 1.645 7.630 1.875 ;
        RECT  4.510 1.645 4.740 2.675 ;
        RECT  4.400 2.335 4.510 2.675 ;
        RECT  2.915 2.405 4.400 2.635 ;
        RECT  3.530 1.745 3.870 2.140 ;
        RECT  1.045 1.745 3.530 1.975 ;
        RECT  2.575 2.365 2.915 2.705 ;
        RECT  0.815 1.345 1.045 3.650 ;
        RECT  0.520 1.345 0.815 1.575 ;
        RECT  0.520 3.420 0.815 3.650 ;
        RECT  0.180 0.940 0.520 1.575 ;
        RECT  0.180 3.420 0.520 3.760 ;
    END
END NOR4BBX4

MACRO NOR4BBX2
    CLASS CORE ;
    FOREIGN NOR4BBX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BBXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.900 0.630 7.130 4.140 ;
        RECT  4.700 0.630 6.900 0.860 ;
        RECT  6.740 3.755 6.900 4.140 ;
        RECT  3.745 3.910 6.740 4.140 ;
        RECT  4.470 0.630 4.700 1.035 ;
        RECT  3.480 0.805 4.470 1.035 ;
        RECT  3.515 3.910 3.745 4.315 ;
        RECT  3.330 3.910 3.515 4.250 ;
        RECT  3.140 0.695 3.480 1.035 ;
        RECT  1.960 0.805 3.140 1.035 ;
        RECT  1.620 0.695 1.960 1.035 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.675 2.395 5.815 2.625 ;
        RECT  5.445 2.395 5.675 3.680 ;
        RECT  1.765 3.450 5.445 3.680 ;
        RECT  1.535 3.450 1.765 3.755 ;
        RECT  1.375 3.450 1.535 3.680 ;
        RECT  1.145 2.340 1.375 3.680 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.005 2.395 5.140 2.625 ;
        RECT  5.005 2.955 5.065 3.195 ;
        RECT  4.835 2.395 5.005 3.195 ;
        RECT  4.775 2.395 4.835 3.185 ;
        RECT  2.160 2.955 4.775 3.185 ;
        RECT  1.875 1.920 2.160 3.185 ;
        RECT  1.820 1.920 1.875 2.260 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.650 1.165 6.460 1.665 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.820 1.265 2.100 ;
        RECT  0.580 1.595 0.905 2.100 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.240 -0.400 7.260 0.400 ;
        RECT  3.900 -0.400 4.240 0.575 ;
        RECT  2.720 -0.400 3.900 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  1.240 -0.400 2.380 0.400 ;
        RECT  0.900 -0.400 1.240 0.895 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.110 4.640 7.260 5.440 ;
        RECT  5.770 4.465 6.110 5.440 ;
        RECT  1.080 4.640 5.770 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.440 1.920 6.670 3.210 ;
        RECT  5.160 1.920 6.440 2.150 ;
        RECT  5.160 1.100 5.420 1.330 ;
        RECT  4.930 1.100 5.160 2.150 ;
        RECT  4.470 1.920 4.930 2.150 ;
        RECT  4.360 1.920 4.470 2.260 ;
        RECT  4.130 1.920 4.360 2.725 ;
        RECT  2.870 2.495 4.130 2.725 ;
        RECT  3.565 1.920 3.675 2.260 ;
        RECT  3.335 1.360 3.565 2.260 ;
        RECT  1.385 1.360 3.335 1.590 ;
        RECT  2.640 1.920 2.870 2.725 ;
        RECT  2.530 1.920 2.640 2.260 ;
        RECT  1.155 1.130 1.385 1.590 ;
        RECT  0.520 1.130 1.155 1.360 ;
        RECT  0.350 0.910 0.520 1.360 ;
        RECT  0.350 2.870 0.520 3.680 ;
        RECT  0.120 0.910 0.350 3.680 ;
    END
END NOR4BBX2

MACRO NOR4BBX1
    CLASS CORE ;
    FOREIGN NOR4BBX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BBXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.930 0.805 5.160 3.755 ;
        RECT  3.350 0.805 4.930 1.035 ;
        RECT  3.825 3.525 4.930 3.755 ;
        RECT  3.485 3.525 3.825 3.865 ;
        RECT  3.065 0.805 3.350 1.425 ;
        RECT  3.010 0.935 3.065 1.425 ;
        RECT  1.575 0.935 3.010 1.275 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.520 2.405 1.765 2.635 ;
        RECT  1.290 1.650 1.520 2.635 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 2.405 2.425 2.635 ;
        RECT  2.110 1.730 2.340 2.635 ;
        RECT  1.905 1.730 2.110 2.070 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 2.275 4.205 2.615 ;
        RECT  3.855 2.275 4.085 3.195 ;
        RECT  3.515 2.940 3.855 3.195 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.175 1.840 0.515 2.500 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 -0.400 5.280 0.400 ;
        RECT  3.770 -0.400 4.110 0.575 ;
        RECT  2.770 -0.400 3.770 0.400 ;
        RECT  2.430 -0.400 2.770 0.575 ;
        RECT  1.155 -0.400 2.430 0.400 ;
        RECT  0.815 -0.400 1.155 0.575 ;
        RECT  0.000 -0.400 0.815 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.715 4.640 5.280 5.440 ;
        RECT  4.375 4.015 4.715 5.440 ;
        RECT  1.265 4.640 4.375 5.440 ;
        RECT  0.925 4.410 1.265 5.440 ;
        RECT  0.000 4.640 0.925 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.455 1.265 4.685 3.190 ;
        RECT  2.915 1.780 4.455 2.010 ;
        RECT  4.315 2.850 4.455 3.190 ;
        RECT  3.245 2.275 3.585 2.620 ;
        RECT  3.005 2.390 3.245 2.620 ;
        RECT  2.775 2.390 3.005 3.125 ;
        RECT  2.575 1.780 2.915 2.160 ;
        RECT  0.990 2.895 2.775 3.125 ;
        RECT  0.760 1.225 0.990 3.125 ;
        RECT  0.520 1.225 0.760 1.455 ;
        RECT  0.520 2.810 0.760 3.125 ;
        RECT  0.180 1.115 0.520 1.455 ;
        RECT  0.180 2.810 0.520 3.150 ;
    END
END NOR4BBX1

MACRO NOR4BXL
    CLASS CORE ;
    FOREIGN NOR4BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.730 1.845 3.745 2.075 ;
        RECT  3.500 1.205 3.730 3.365 ;
        RECT  3.200 1.205 3.500 1.435 ;
        RECT  3.300 3.025 3.500 3.365 ;
        RECT  1.540 1.095 3.200 1.435 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 2.335 1.440 3.170 ;
        RECT  1.105 2.940 1.210 3.170 ;
        RECT  0.875 2.940 1.105 3.195 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 2.340 2.170 2.680 ;
        RECT  1.830 1.845 1.900 2.680 ;
        RECT  1.670 1.845 1.830 2.570 ;
        RECT  1.535 1.845 1.670 2.075 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 1.735 3.160 2.155 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.135 1.660 0.520 2.235 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 -0.400 3.960 0.400 ;
        RECT  3.420 -0.400 3.760 0.575 ;
        RECT  2.440 -0.400 3.420 0.400 ;
        RECT  2.100 -0.400 2.440 0.575 ;
        RECT  1.180 -0.400 2.100 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 4.640 3.960 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.630 2.495 3.270 2.725 ;
        RECT  2.400 2.495 2.630 3.680 ;
        RECT  0.520 3.450 2.400 3.680 ;
        RECT  0.750 1.145 0.980 2.700 ;
        RECT  0.520 1.145 0.750 1.375 ;
        RECT  0.520 2.470 0.750 2.700 ;
        RECT  0.180 1.025 0.520 1.375 ;
        RECT  0.290 2.470 0.520 3.680 ;
        RECT  0.180 3.025 0.290 3.365 ;
    END
END NOR4BXL

MACRO NOR4BX4
    CLASS CORE ;
    FOREIGN NOR4BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 2.380 11.740 3.780 ;
        RECT  11.435 1.185 11.665 3.875 ;
        RECT  10.795 1.185 11.435 1.415 ;
        RECT  11.360 2.380 11.435 3.875 ;
        RECT  8.885 3.645 11.360 3.875 ;
        RECT  10.455 1.075 10.795 1.415 ;
        RECT  9.340 1.185 10.455 1.415 ;
        RECT  9.000 1.075 9.340 1.415 ;
        RECT  3.400 1.185 9.000 1.415 ;
        RECT  8.775 3.640 8.885 3.980 ;
        RECT  8.545 3.640 8.775 4.235 ;
        RECT  3.825 4.005 8.545 4.235 ;
        RECT  3.485 4.005 3.825 4.345 ;
        RECT  3.060 1.075 3.400 1.415 ;
        RECT  1.960 1.185 3.060 1.415 ;
        RECT  1.620 1.075 1.960 1.415 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.025 1.800 11.165 2.140 ;
        RECT  10.795 1.800 11.025 3.185 ;
        RECT  6.385 2.955 10.795 3.185 ;
        RECT  6.330 2.955 6.385 3.195 ;
        RECT  6.220 2.595 6.330 3.195 ;
        RECT  5.990 2.595 6.220 3.775 ;
        RECT  1.520 3.545 5.990 3.775 ;
        RECT  1.290 2.210 1.520 3.775 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.355 2.000 10.465 2.405 ;
        RECT  10.125 2.000 10.355 2.720 ;
        RECT  7.220 2.490 10.125 2.720 ;
        RECT  6.990 2.110 7.220 2.720 ;
        RECT  6.880 2.110 6.990 2.450 ;
        RECT  6.740 2.110 6.880 2.405 ;
        RECT  5.490 2.110 6.740 2.340 ;
        RECT  5.380 2.110 5.490 2.450 ;
        RECT  5.140 2.110 5.380 3.315 ;
        RECT  4.835 2.965 5.140 3.315 ;
        RECT  2.245 3.085 4.835 3.315 ;
        RECT  1.960 2.335 2.245 3.315 ;
        RECT  1.905 2.335 1.960 2.675 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 1.920 9.795 2.260 ;
        RECT  8.135 2.030 9.455 2.260 ;
        RECT  7.860 1.820 8.135 2.260 ;
        RECT  7.630 1.645 7.860 2.260 ;
        RECT  4.740 1.645 7.630 1.875 ;
        RECT  4.510 1.645 4.740 2.675 ;
        RECT  4.400 2.335 4.510 2.675 ;
        RECT  2.915 2.405 4.400 2.635 ;
        RECT  2.575 2.365 2.915 2.705 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.170 1.845 0.510 2.555 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.530 -0.400 11.880 0.400 ;
        RECT  11.190 -0.400 11.530 0.955 ;
        RECT  10.065 -0.400 11.190 0.400 ;
        RECT  9.725 -0.400 10.065 0.955 ;
        RECT  8.620 -0.400 9.725 0.400 ;
        RECT  8.280 -0.400 8.620 0.955 ;
        RECT  4.135 -0.400 8.280 0.400 ;
        RECT  3.795 -0.400 4.135 0.955 ;
        RECT  2.680 -0.400 3.795 0.400 ;
        RECT  2.340 -0.400 2.680 0.950 ;
        RECT  1.240 -0.400 2.340 0.400 ;
        RECT  0.900 -0.400 1.240 0.950 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.530 4.640 11.880 5.440 ;
        RECT  11.190 4.465 11.530 5.440 ;
        RECT  6.355 4.640 11.190 5.440 ;
        RECT  6.015 4.465 6.355 5.440 ;
        RECT  1.295 4.640 6.015 5.440 ;
        RECT  0.955 4.465 1.295 5.440 ;
        RECT  0.000 4.640 0.955 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.530 1.745 3.870 2.140 ;
        RECT  1.045 1.745 3.530 1.975 ;
        RECT  0.815 1.345 1.045 3.650 ;
        RECT  0.520 1.345 0.815 1.575 ;
        RECT  0.520 3.420 0.815 3.650 ;
        RECT  0.180 0.940 0.520 1.575 ;
        RECT  0.180 3.420 0.520 3.760 ;
    END
END NOR4BX4

MACRO NOR4BX2
    CLASS CORE ;
    FOREIGN NOR4BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.140 0.805 6.370 3.755 ;
        RECT  6.080 0.805 6.140 1.285 ;
        RECT  4.180 3.525 6.140 3.755 ;
        RECT  3.480 0.805 6.080 1.035 ;
        RECT  3.880 3.500 4.180 3.780 ;
        RECT  3.540 3.470 3.880 3.810 ;
        RECT  3.140 0.750 3.480 1.090 ;
        RECT  1.620 0.805 3.140 1.035 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.795 2.340 5.910 2.680 ;
        RECT  5.570 2.340 5.795 3.195 ;
        RECT  5.565 2.395 5.570 3.195 ;
        RECT  1.535 2.965 5.565 3.195 ;
        RECT  1.430 2.940 1.535 3.195 ;
        RECT  1.090 2.390 1.430 3.195 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.425 1.665 5.725 2.100 ;
        RECT  5.135 1.440 5.425 2.100 ;
        RECT  2.500 1.440 5.135 1.670 ;
        RECT  2.350 1.440 2.500 1.845 ;
        RECT  2.120 1.440 2.350 2.240 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.900 4.680 2.635 ;
        RECT  3.080 1.900 4.175 2.130 ;
        RECT  2.740 1.900 3.080 2.240 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.815 1.820 1.180 2.155 ;
        RECT  0.585 1.660 0.815 2.155 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.240 -0.400 6.600 0.400 ;
        RECT  3.900 -0.400 4.240 0.575 ;
        RECT  2.720 -0.400 3.900 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  1.240 -0.400 2.380 0.400 ;
        RECT  0.900 -0.400 1.240 0.895 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 4.640 6.600 5.440 ;
        RECT  5.980 4.465 6.320 5.440 ;
        RECT  1.200 4.640 5.980 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.395 2.395 3.750 2.700 ;
        RECT  1.890 2.470 3.395 2.700 ;
        RECT  1.660 1.265 1.890 2.700 ;
        RECT  1.315 1.265 1.660 1.495 ;
        RECT  1.085 1.125 1.315 1.495 ;
        RECT  0.520 1.125 1.085 1.355 ;
        RECT  0.355 0.910 0.520 1.355 ;
        RECT  0.355 2.870 0.520 3.680 ;
        RECT  0.125 0.910 0.355 3.680 ;
    END
END NOR4BX2

MACRO NOR4BX1
    CLASS CORE ;
    FOREIGN NOR4BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.730 1.845 3.745 2.075 ;
        RECT  3.500 1.210 3.730 3.355 ;
        RECT  3.200 1.210 3.500 1.440 ;
        RECT  3.300 3.015 3.500 3.355 ;
        RECT  1.540 1.100 3.200 1.440 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 2.335 1.440 3.170 ;
        RECT  1.105 2.940 1.210 3.170 ;
        RECT  0.875 2.940 1.105 3.195 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 2.340 2.170 2.680 ;
        RECT  1.830 1.845 1.900 2.680 ;
        RECT  1.670 1.845 1.830 2.570 ;
        RECT  1.535 1.845 1.670 2.075 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 1.735 3.160 2.155 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.515 1.660 0.520 2.230 ;
        RECT  0.175 1.660 0.515 2.235 ;
        RECT  0.135 1.660 0.175 2.230 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 -0.400 3.960 0.400 ;
        RECT  3.420 -0.400 3.760 0.575 ;
        RECT  2.440 -0.400 3.420 0.400 ;
        RECT  2.100 -0.400 2.440 0.575 ;
        RECT  1.180 -0.400 2.100 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 3.960 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.630 2.495 3.270 2.725 ;
        RECT  2.400 2.495 2.630 3.680 ;
        RECT  0.520 3.450 2.400 3.680 ;
        RECT  0.750 1.145 0.980 2.700 ;
        RECT  0.520 1.145 0.750 1.375 ;
        RECT  0.520 2.470 0.750 2.700 ;
        RECT  0.180 1.035 0.520 1.375 ;
        RECT  0.290 2.470 0.520 3.680 ;
        RECT  0.180 2.970 0.290 3.310 ;
    END
END NOR4BX1

MACRO NOR4XL
    CLASS CORE ;
    FOREIGN NOR4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.130 3.745 3.195 ;
        RECT  0.940 1.130 3.515 1.470 ;
        RECT  3.165 2.965 3.515 3.195 ;
        RECT  2.825 2.930 3.165 3.740 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.310 0.570 2.975 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.770 1.585 2.210 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 1.820 2.325 2.160 ;
        RECT  1.905 1.820 2.135 3.195 ;
        RECT  1.535 2.940 1.905 3.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 2.075 3.260 2.590 ;
        RECT  2.920 1.845 3.160 2.590 ;
        RECT  2.855 1.845 2.920 2.075 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 3.960 0.400 ;
        RECT  3.440 -0.400 3.780 0.575 ;
        RECT  2.200 -0.400 3.440 0.400 ;
        RECT  1.860 -0.400 2.200 0.575 ;
        RECT  0.520 -0.400 1.860 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 3.960 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR4XL

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4XL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.005 2.380 11.080 3.780 ;
        RECT  10.775 1.185 11.005 3.875 ;
        RECT  10.135 1.185 10.775 1.415 ;
        RECT  10.700 2.380 10.775 3.875 ;
        RECT  8.225 3.645 10.700 3.875 ;
        RECT  9.795 1.075 10.135 1.415 ;
        RECT  8.680 1.185 9.795 1.415 ;
        RECT  8.340 1.075 8.680 1.415 ;
        RECT  2.725 1.185 8.340 1.415 ;
        RECT  8.115 3.640 8.225 3.980 ;
        RECT  7.885 3.640 8.115 4.235 ;
        RECT  3.165 4.005 7.885 4.235 ;
        RECT  2.825 4.005 3.165 4.345 ;
        RECT  2.385 1.075 2.725 1.415 ;
        RECT  1.255 1.185 2.385 1.415 ;
        RECT  0.915 1.075 1.255 1.415 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.365 1.800 10.505 2.140 ;
        RECT  10.135 1.800 10.365 3.185 ;
        RECT  5.670 2.955 10.135 3.185 ;
        RECT  5.560 2.595 5.670 3.185 ;
        RECT  5.330 2.595 5.560 3.775 ;
        RECT  0.885 3.545 5.330 3.775 ;
        RECT  0.655 2.335 0.885 3.775 ;
        RECT  0.205 2.335 0.655 2.675 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.695 2.000 9.805 2.405 ;
        RECT  9.465 2.000 9.695 2.720 ;
        RECT  6.560 2.490 9.465 2.720 ;
        RECT  6.330 2.110 6.560 2.720 ;
        RECT  6.080 2.110 6.330 2.450 ;
        RECT  4.830 2.110 6.080 2.340 ;
        RECT  4.720 2.110 4.830 2.450 ;
        RECT  4.490 2.110 4.720 3.315 ;
        RECT  4.405 2.940 4.490 3.315 ;
        RECT  1.765 3.085 4.405 3.315 ;
        RECT  1.585 2.965 1.765 3.315 ;
        RECT  1.355 2.335 1.585 3.315 ;
        RECT  1.245 2.335 1.355 2.675 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.795 1.920 9.135 2.260 ;
        RECT  7.475 2.030 8.795 2.260 ;
        RECT  7.200 1.820 7.475 2.260 ;
        RECT  6.970 1.645 7.200 2.260 ;
        RECT  4.080 1.645 6.970 1.875 ;
        RECT  3.740 1.645 4.080 2.675 ;
        RECT  2.425 1.645 3.740 1.875 ;
        RECT  2.255 1.645 2.425 2.075 ;
        RECT  1.915 1.645 2.255 2.260 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 2.405 3.210 2.850 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.870 -0.400 11.220 0.400 ;
        RECT  10.530 -0.400 10.870 0.955 ;
        RECT  9.405 -0.400 10.530 0.400 ;
        RECT  9.065 -0.400 9.405 0.955 ;
        RECT  7.960 -0.400 9.065 0.400 ;
        RECT  7.620 -0.400 7.960 0.955 ;
        RECT  3.460 -0.400 7.620 0.400 ;
        RECT  3.120 -0.400 3.460 0.955 ;
        RECT  1.985 -0.400 3.120 0.400 ;
        RECT  1.645 -0.400 1.985 0.950 ;
        RECT  0.520 -0.400 1.645 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.870 4.640 11.220 5.440 ;
        RECT  10.530 4.465 10.870 5.440 ;
        RECT  5.695 4.640 10.530 5.440 ;
        RECT  5.355 4.465 5.695 5.440 ;
        RECT  0.520 4.640 5.355 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.205 5.725 4.235 ;
        RECT  3.020 1.205 5.495 1.435 ;
        RECT  5.420 3.755 5.495 4.235 ;
        RECT  3.165 4.005 5.420 4.235 ;
        RECT  2.825 4.005 3.165 4.345 ;
        RECT  2.680 1.095 3.020 1.435 ;
        RECT  1.255 1.205 2.680 1.435 ;
        RECT  0.915 1.095 1.255 1.435 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 2.335 5.260 2.675 ;
        RECT  4.920 2.335 5.150 3.775 ;
        RECT  0.885 3.545 4.920 3.775 ;
        RECT  0.655 2.335 0.885 3.775 ;
        RECT  0.205 2.335 0.655 2.675 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.360 1.665 4.590 3.315 ;
        RECT  4.250 1.665 4.360 2.005 ;
        RECT  1.765 3.085 4.360 3.315 ;
        RECT  1.585 2.965 1.765 3.315 ;
        RECT  1.355 2.335 1.585 3.315 ;
        RECT  1.245 2.335 1.355 2.675 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 2.335 4.080 2.675 ;
        RECT  3.740 1.865 3.970 2.675 ;
        RECT  2.425 1.865 3.740 2.095 ;
        RECT  2.255 1.845 2.425 2.095 ;
        RECT  1.920 1.845 2.255 2.260 ;
        RECT  1.915 1.920 1.920 2.260 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 2.330 3.260 2.670 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 5.940 0.400 ;
        RECT  3.440 -0.400 3.780 0.575 ;
        RECT  2.200 -0.400 3.440 0.400 ;
        RECT  1.860 -0.400 2.200 0.575 ;
        RECT  0.520 -0.400 1.860 0.400 ;
        RECT  0.180 -0.400 0.520 1.010 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.695 4.640 5.940 5.440 ;
        RECT  5.355 4.465 5.695 5.440 ;
        RECT  0.520 4.640 5.355 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR4X2

MACRO NOR4X1
    CLASS CORE ;
    FOREIGN NOR4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.130 3.745 3.195 ;
        RECT  0.940 1.130 3.515 1.470 ;
        RECT  3.165 2.965 3.515 3.195 ;
        RECT  2.825 2.930 3.165 3.740 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 2.275 0.565 2.615 ;
        RECT  0.225 2.275 0.560 2.940 ;
        RECT  0.205 2.405 0.225 2.635 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.770 1.585 2.180 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 1.820 2.255 2.160 ;
        RECT  1.905 1.820 2.135 3.195 ;
        RECT  1.535 2.940 1.905 3.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 1.765 3.260 2.350 ;
        RECT  2.855 1.845 2.920 2.075 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 3.960 0.400 ;
        RECT  3.440 -0.400 3.780 0.575 ;
        RECT  2.200 -0.400 3.440 0.400 ;
        RECT  1.860 -0.400 2.200 0.575 ;
        RECT  0.520 -0.400 1.860 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 3.960 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR4X1

MACRO NOR3BXL
    CLASS CORE ;
    FOREIGN NOR3BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 1.130 3.780 3.755 ;
        RECT  1.750 1.130 3.550 1.470 ;
        RECT  3.515 3.195 3.550 3.755 ;
        RECT  3.440 3.195 3.515 3.690 ;
        RECT  2.820 3.350 3.440 3.690 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.760 2.405 1.765 2.635 ;
        RECT  1.105 2.250 1.760 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.740 2.720 2.145 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 1.285 1.105 1.515 ;
        RECT  0.800 1.285 1.030 1.920 ;
        RECT  0.655 1.580 0.800 1.920 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 -0.400 3.960 0.400 ;
        RECT  2.510 -0.400 2.850 0.575 ;
        RECT  1.495 -0.400 2.510 0.400 ;
        RECT  1.155 -0.400 1.495 0.575 ;
        RECT  0.000 -0.400 1.155 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 4.640 3.960 5.440 ;
        RECT  0.960 3.350 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 2.250 3.300 2.590 ;
        RECT  2.960 2.250 3.190 3.120 ;
        RECT  0.520 2.890 2.960 3.120 ;
        RECT  0.410 0.995 0.540 1.350 ;
        RECT  0.410 2.790 0.520 3.130 ;
        RECT  0.180 0.995 0.410 3.130 ;
    END
END NOR3BXL

MACRO NOR3BX4
    CLASS CORE ;
    FOREIGN NOR3BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3BXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.970 1.820 7.120 3.580 ;
        RECT  6.740 1.125 6.970 3.580 ;
        RECT  5.195 1.125 6.740 1.355 ;
        RECT  6.560 3.240 6.740 3.580 ;
        RECT  3.820 3.240 6.560 3.470 ;
        RECT  4.965 0.695 5.195 1.355 ;
        RECT  4.855 0.695 4.965 1.035 ;
        RECT  3.670 0.805 4.855 1.035 ;
        RECT  3.745 3.240 3.820 3.525 ;
        RECT  3.515 3.240 3.745 3.640 ;
        RECT  3.330 0.695 3.670 1.035 ;
        RECT  3.180 3.410 3.515 3.640 ;
        RECT  2.150 0.805 3.330 1.035 ;
        RECT  2.840 3.410 3.180 3.750 ;
        RECT  1.810 0.695 2.150 1.035 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.700 1.740 5.280 2.080 ;
        RECT  4.470 1.265 4.700 2.080 ;
        RECT  1.765 1.265 4.470 1.495 ;
        RECT  1.535 1.265 1.765 2.635 ;
        RECT  1.330 2.250 1.535 2.590 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.665 2.195 5.895 2.545 ;
        RECT  4.095 2.315 5.665 2.545 ;
        RECT  3.985 2.185 4.095 2.545 ;
        RECT  3.755 1.725 3.985 2.545 ;
        RECT  3.745 1.725 3.755 2.100 ;
        RECT  2.425 1.725 3.745 1.955 ;
        RECT  2.390 1.725 2.425 2.155 ;
        RECT  2.050 1.725 2.390 2.160 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 1.285 1.105 1.515 ;
        RECT  0.800 1.285 1.030 2.180 ;
        RECT  0.655 1.840 0.800 2.180 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.915 -0.400 7.260 0.400 ;
        RECT  5.575 -0.400 5.915 0.895 ;
        RECT  4.435 -0.400 5.575 0.400 ;
        RECT  4.095 -0.400 4.435 0.575 ;
        RECT  2.910 -0.400 4.095 0.400 ;
        RECT  2.570 -0.400 2.910 0.575 ;
        RECT  1.430 -0.400 2.570 0.400 ;
        RECT  1.090 -0.400 1.430 0.895 ;
        RECT  0.000 -0.400 1.090 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.040 4.640 7.260 5.440 ;
        RECT  4.700 3.765 5.040 5.440 ;
        RECT  1.300 4.640 4.700 5.440 ;
        RECT  0.960 3.575 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.125 1.585 6.420 3.005 ;
        RECT  6.050 1.585 6.125 1.835 ;
        RECT  3.190 2.775 6.125 3.005 ;
        RECT  2.830 2.185 3.190 3.175 ;
        RECT  0.520 2.945 2.830 3.175 ;
        RECT  0.410 0.830 0.570 1.185 ;
        RECT  0.410 2.945 0.520 3.320 ;
        RECT  0.180 0.830 0.410 3.320 ;
    END
END NOR3BX4

MACRO NOR3BX2
    CLASS CORE ;
    FOREIGN NOR3BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.790 0.805 5.020 3.615 ;
        RECT  4.760 0.805 4.790 1.285 ;
        RECT  4.760 3.195 4.790 3.615 ;
        RECT  3.670 0.805 4.760 1.035 ;
        RECT  3.745 3.385 4.760 3.615 ;
        RECT  3.515 3.385 3.745 3.755 ;
        RECT  3.330 0.695 3.670 1.035 ;
        RECT  3.180 3.385 3.515 3.615 ;
        RECT  2.150 0.805 3.330 1.035 ;
        RECT  2.840 3.385 3.180 3.760 ;
        RECT  1.810 0.695 2.150 1.035 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.655 4.560 1.995 ;
        RECT  4.220 1.360 4.450 1.995 ;
        RECT  1.760 1.360 4.220 1.590 ;
        RECT  1.760 2.405 1.765 2.635 ;
        RECT  1.530 1.360 1.760 2.635 ;
        RECT  1.460 2.075 1.530 2.635 ;
        RECT  1.375 2.250 1.460 2.635 ;
        RECT  1.265 2.250 1.375 2.590 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 2.330 4.095 2.670 ;
        RECT  3.755 1.935 3.985 2.670 ;
        RECT  2.425 1.935 3.755 2.165 ;
        RECT  2.335 1.845 2.425 2.165 ;
        RECT  2.105 1.845 2.335 2.275 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 1.285 1.105 1.515 ;
        RECT  0.800 1.285 1.030 1.920 ;
        RECT  0.655 1.580 0.800 1.920 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 -0.400 5.280 0.400 ;
        RECT  2.570 -0.400 2.910 0.575 ;
        RECT  1.430 -0.400 2.570 0.400 ;
        RECT  1.090 -0.400 1.430 0.895 ;
        RECT  0.000 -0.400 1.090 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.040 4.640 5.280 5.440 ;
        RECT  4.700 3.850 5.040 5.440 ;
        RECT  1.300 4.640 4.700 5.440 ;
        RECT  0.960 3.705 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 2.395 3.300 2.625 ;
        RECT  2.960 2.395 3.190 3.155 ;
        RECT  0.520 2.925 2.960 3.155 ;
        RECT  0.410 0.830 0.570 1.185 ;
        RECT  0.410 2.815 0.520 3.155 ;
        RECT  0.180 0.830 0.410 3.155 ;
    END
END NOR3BX2

MACRO NOR3BX1
    CLASS CORE ;
    FOREIGN NOR3BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.610 1.130 3.840 3.755 ;
        RECT  1.750 1.130 3.610 1.470 ;
        RECT  3.160 3.525 3.610 3.755 ;
        RECT  2.820 3.525 3.160 3.880 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.760 2.405 1.765 2.635 ;
        RECT  1.105 2.250 1.760 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.740 2.720 2.145 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 1.285 1.105 1.515 ;
        RECT  0.800 1.285 1.030 1.920 ;
        RECT  0.655 1.580 0.800 1.920 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 -0.400 3.960 0.400 ;
        RECT  2.510 -0.400 2.850 0.575 ;
        RECT  1.495 -0.400 2.510 0.400 ;
        RECT  1.155 -0.400 1.495 0.575 ;
        RECT  0.000 -0.400 1.155 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 4.640 3.960 5.440 ;
        RECT  0.960 3.705 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 2.250 3.300 2.590 ;
        RECT  2.960 2.250 3.190 3.155 ;
        RECT  0.520 2.925 2.960 3.155 ;
        RECT  0.410 0.995 0.540 1.350 ;
        RECT  0.410 2.815 0.520 3.155 ;
        RECT  0.180 0.995 0.410 3.155 ;
    END
END NOR3BX1

MACRO NOR3XL
    CLASS CORE ;
    FOREIGN NOR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 1.185 2.520 3.755 ;
        RECT  2.290 1.185 2.510 3.835 ;
        RECT  0.740 1.185 2.290 1.525 ;
        RECT  2.100 3.480 2.290 3.835 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.180 2.405 0.520 3.070 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.770 1.360 2.355 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 2.305 2.060 2.645 ;
        RECT  1.720 2.305 1.950 3.195 ;
        RECT  1.535 2.965 1.720 3.195 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 2.640 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 2.640 5.440 ;
        RECT  0.180 3.505 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR3XL

MACRO NOR3X4
    CLASS CORE ;
    FOREIGN NOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 2.380 6.460 3.780 ;
        RECT  6.080 1.125 6.310 3.780 ;
        RECT  4.120 1.125 6.080 1.355 ;
        RECT  5.725 3.400 6.080 3.745 ;
        RECT  2.440 3.515 5.725 3.745 ;
        RECT  3.780 1.015 4.120 1.355 ;
        RECT  2.680 1.125 3.780 1.355 ;
        RECT  2.340 1.015 2.680 1.355 ;
        RECT  2.100 3.515 2.440 3.855 ;
        RECT  1.240 1.125 2.340 1.355 ;
        RECT  0.900 1.015 1.240 1.355 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 2.510 4.360 3.250 ;
        RECT  3.745 2.940 4.005 3.250 ;
        RECT  0.560 3.020 3.745 3.250 ;
        RECT  0.330 2.210 0.560 3.250 ;
        RECT  0.205 2.210 0.330 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.560 2.050 5.095 2.280 ;
        RECT  3.330 2.050 3.560 2.560 ;
        RECT  1.480 2.330 3.330 2.560 ;
        RECT  1.370 2.130 1.480 2.560 ;
        RECT  1.140 1.845 1.370 2.560 ;
        RECT  0.875 1.845 1.140 2.075 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.695 2.440 5.800 2.780 ;
        RECT  5.465 1.590 5.695 2.780 ;
        RECT  2.680 1.590 5.465 1.820 ;
        RECT  5.460 2.440 5.465 2.780 ;
        RECT  2.340 1.590 2.680 2.085 ;
        RECT  2.195 1.800 2.340 2.075 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.840 -0.400 6.600 0.400 ;
        RECT  4.500 -0.400 4.840 0.895 ;
        RECT  3.400 -0.400 4.500 0.400 ;
        RECT  3.060 -0.400 3.400 0.895 ;
        RECT  1.960 -0.400 3.060 0.400 ;
        RECT  1.620 -0.400 1.960 0.895 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 4.640 6.600 5.440 ;
        RECT  3.990 4.090 4.330 5.440 ;
        RECT  0.520 4.640 3.990 5.440 ;
        RECT  0.180 3.840 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR3X4

MACRO NOR3X2
    CLASS CORE ;
    FOREIGN NOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.070 4.405 3.590 ;
        RECT  2.680 1.070 4.175 1.300 ;
        RECT  4.100 3.220 4.175 3.590 ;
        RECT  2.440 3.360 4.100 3.590 ;
        RECT  2.340 0.635 2.680 1.445 ;
        RECT  2.100 3.360 2.440 3.740 ;
        RECT  1.240 1.215 2.340 1.445 ;
        RECT  0.900 0.635 1.240 1.445 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 2.255 3.865 3.125 ;
        RECT  0.760 2.895 3.580 3.125 ;
        RECT  0.530 2.405 0.760 3.125 ;
        RECT  0.420 2.405 0.530 2.970 ;
        RECT  0.205 2.405 0.420 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.245 1.585 3.350 1.925 ;
        RECT  3.015 1.585 3.245 2.665 ;
        RECT  3.010 1.585 3.015 1.925 ;
        RECT  1.480 2.435 3.015 2.665 ;
        RECT  1.475 1.925 1.480 2.665 ;
        RECT  1.250 1.870 1.475 2.665 ;
        RECT  1.140 1.870 1.250 2.265 ;
        RECT  1.105 1.870 1.140 2.100 ;
        RECT  0.875 1.845 1.105 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.845 2.425 2.205 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 -0.400 4.620 0.400 ;
        RECT  1.620 -0.400 1.960 0.950 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 4.640 4.620 5.440 ;
        RECT  3.940 3.820 4.280 5.440 ;
        RECT  0.520 4.640 3.940 5.440 ;
        RECT  0.180 3.615 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR3X2

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 1.130 2.520 3.755 ;
        RECT  2.290 1.130 2.510 3.880 ;
        RECT  0.740 1.130 2.290 1.470 ;
        RECT  2.100 3.525 2.290 3.880 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.515 2.250 0.520 2.590 ;
        RECT  0.180 2.250 0.515 2.915 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.770 1.360 2.355 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 2.250 2.060 2.590 ;
        RECT  1.720 2.250 1.950 3.195 ;
        RECT  1.535 2.965 1.720 3.195 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 2.640 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.520 -0.400 1.300 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 2.640 5.440 ;
        RECT  0.180 3.715 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR3X1

MACRO NOR2BXL
    CLASS CORE ;
    FOREIGN NOR2BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.280 1.240 2.510 3.350 ;
        RECT  1.890 1.240 2.280 1.470 ;
        RECT  2.120 2.965 2.280 3.350 ;
        RECT  1.550 1.130 1.890 1.470 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.550 2.380 1.980 2.660 ;
        RECT  1.210 2.380 1.550 2.780 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.520 2.440 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 -0.400 2.640 0.400 ;
        RECT  2.120 -0.400 2.460 0.575 ;
        RECT  1.180 -0.400 2.120 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.140 4.640 2.640 5.440 ;
        RECT  0.800 4.465 1.140 5.440 ;
        RECT  0.000 4.640 0.800 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.980 1.770 2.050 2.110 ;
        RECT  0.750 1.350 0.980 3.200 ;
        RECT  0.520 1.350 0.750 1.580 ;
        RECT  0.520 2.970 0.750 3.200 ;
        RECT  0.180 1.240 0.520 1.580 ;
        RECT  0.180 2.970 0.520 3.310 ;
    END
END NOR2BXL

MACRO NOR2BX4
    CLASS CORE ;
    FOREIGN NOR2BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.760 1.110 5.140 3.300 ;
        RECT  3.670 1.110 4.760 1.410 ;
        RECT  4.720 2.910 4.760 3.300 ;
        RECT  2.160 2.960 4.720 3.300 ;
        RECT  3.330 1.070 3.670 1.410 ;
        RECT  2.150 1.180 3.330 1.410 ;
        RECT  1.810 1.070 2.150 1.410 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 2.365 3.870 2.730 ;
        RECT  1.765 2.500 3.530 2.730 ;
        RECT  1.550 2.375 1.765 2.730 ;
        RECT  1.210 2.190 1.550 2.730 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 1.830 0.520 2.400 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 -0.400 5.280 0.400 ;
        RECT  4.100 -0.400 4.440 0.575 ;
        RECT  2.910 -0.400 4.100 0.400 ;
        RECT  2.570 -0.400 2.910 0.575 ;
        RECT  1.380 -0.400 2.570 0.400 ;
        RECT  1.040 -0.400 1.380 0.575 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 4.640 5.280 5.440 ;
        RECT  3.480 4.465 3.820 5.440 ;
        RECT  1.180 4.630 3.480 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.295 1.645 4.525 2.295 ;
        RECT  2.520 1.645 4.295 1.875 ;
        RECT  2.180 1.645 2.520 2.260 ;
        RECT  0.980 1.645 2.180 1.875 ;
        RECT  0.750 1.290 0.980 3.560 ;
        RECT  0.620 1.290 0.750 1.520 ;
        RECT  0.520 3.330 0.750 3.560 ;
        RECT  0.280 1.180 0.620 1.520 ;
        RECT  0.180 3.330 0.520 3.670 ;
    END
END NOR2BX4

MACRO NOR2BX2
    CLASS CORE ;
    FOREIGN NOR2BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.295 3.820 3.220 ;
        RECT  3.060 1.295 3.590 1.525 ;
        RECT  3.515 2.965 3.590 3.220 ;
        RECT  2.480 2.990 3.515 3.220 ;
        RECT  2.720 1.185 3.060 1.525 ;
        RECT  2.140 2.990 2.480 3.330 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.050 1.755 3.340 2.375 ;
        RECT  1.840 1.755 3.050 1.985 ;
        RECT  1.570 1.260 1.840 1.985 ;
        RECT  1.460 1.260 1.570 2.160 ;
        RECT  1.285 1.755 1.460 2.160 ;
        RECT  1.230 1.820 1.285 2.160 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.180 1.920 0.520 2.660 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 3.960 0.400 ;
        RECT  3.440 -0.400 3.780 1.020 ;
        RECT  2.290 -0.400 3.440 0.400 ;
        RECT  1.950 -0.400 2.290 0.575 ;
        RECT  0.000 -0.400 1.950 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 4.640 3.960 5.440 ;
        RECT  3.440 4.465 3.780 5.440 ;
        RECT  1.160 4.640 3.440 5.440 ;
        RECT  0.820 4.465 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.240 2.260 2.580 2.630 ;
        RECT  0.980 2.400 2.240 2.630 ;
        RECT  0.750 1.310 0.980 3.370 ;
        RECT  0.520 1.310 0.750 1.540 ;
        RECT  0.520 3.140 0.750 3.370 ;
        RECT  0.180 1.200 0.520 1.540 ;
        RECT  0.180 3.140 0.520 3.480 ;
    END
END NOR2BX2

MACRO NOR2BX1
    CLASS CORE ;
    FOREIGN NOR2BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2BXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.280 1.240 2.510 3.605 ;
        RECT  1.890 1.240 2.280 1.470 ;
        RECT  2.120 2.965 2.280 3.605 ;
        RECT  1.550 1.130 1.890 1.470 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.550 2.380 1.980 2.660 ;
        RECT  1.210 2.380 1.550 2.815 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.040 0.520 2.660 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 -0.400 2.640 0.400 ;
        RECT  2.120 -0.400 2.460 0.575 ;
        RECT  1.330 -0.400 2.120 0.400 ;
        RECT  0.990 -0.400 1.330 0.575 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.140 4.640 2.640 5.440 ;
        RECT  0.800 3.785 1.140 5.440 ;
        RECT  0.000 4.640 0.800 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.740 1.805 2.050 2.145 ;
        RECT  0.980 1.860 1.740 2.090 ;
        RECT  0.750 1.355 0.980 3.235 ;
        RECT  0.520 1.355 0.750 1.615 ;
        RECT  0.520 3.005 0.750 3.235 ;
        RECT  0.180 1.275 0.520 1.615 ;
        RECT  0.180 3.005 0.520 3.345 ;
    END
END NOR2BX1

MACRO NOR2XL
    CLASS CORE ;
    FOREIGN NOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.620 1.240 1.850 3.250 ;
        RECT  1.160 1.240 1.620 1.470 ;
        RECT  1.460 2.630 1.620 3.250 ;
        RECT  0.820 1.130 1.160 1.470 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.380 0.840 2.660 ;
        RECT  0.200 2.300 0.540 2.660 ;
        RECT  0.140 2.380 0.200 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.705 1.390 2.110 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 -0.400 1.980 0.400 ;
        RECT  1.460 -0.400 1.800 0.575 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 1.980 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR2XL

MACRO NOR2X4
    CLASS CORE ;
    FOREIGN NOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.820 4.480 3.220 ;
        RECT  4.420 1.115 4.440 3.220 ;
        RECT  4.140 1.115 4.420 3.530 ;
        RECT  2.720 1.115 4.140 1.415 ;
        RECT  4.100 1.820 4.140 3.530 ;
        RECT  4.080 2.910 4.100 3.530 ;
        RECT  1.520 3.190 4.080 3.530 ;
        RECT  2.380 1.075 2.720 1.415 ;
        RECT  1.280 1.185 2.380 1.415 ;
        RECT  0.940 1.075 1.280 1.415 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 2.355 3.050 2.695 ;
        RECT  2.710 2.355 2.940 2.960 ;
        RECT  1.105 2.730 2.710 2.960 ;
        RECT  0.875 2.730 1.105 3.195 ;
        RECT  0.830 2.730 0.875 2.970 ;
        RECT  0.600 2.065 0.830 2.970 ;
        RECT  0.490 2.065 0.600 2.405 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.750 1.950 3.860 2.290 ;
        RECT  3.520 1.655 3.750 2.290 ;
        RECT  1.860 1.655 3.520 1.885 ;
        RECT  1.630 1.655 1.860 2.205 ;
        RECT  1.535 1.845 1.630 2.205 ;
        RECT  1.520 1.975 1.535 2.205 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.480 -0.400 4.620 0.400 ;
        RECT  3.140 -0.400 3.480 0.575 ;
        RECT  2.000 -0.400 3.140 0.400 ;
        RECT  1.660 -0.400 2.000 0.950 ;
        RECT  0.520 -0.400 1.660 0.400 ;
        RECT  0.180 -0.400 0.520 1.315 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 4.640 4.620 5.440 ;
        RECT  2.840 4.465 3.180 5.440 ;
        RECT  0.540 4.640 2.840 5.440 ;
        RECT  0.200 4.465 0.540 5.440 ;
        RECT  0.000 4.640 0.200 5.440 ;
        END
    END VDD
END NOR2X4

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 1.295 3.180 3.195 ;
        RECT  2.950 1.295 3.160 3.220 ;
        RECT  2.400 1.295 2.950 1.525 ;
        RECT  2.855 2.965 2.950 3.220 ;
        RECT  1.820 2.990 2.855 3.220 ;
        RECT  2.060 0.715 2.400 1.525 ;
        RECT  1.480 2.990 1.820 3.330 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.390 1.755 2.720 2.370 ;
        RECT  0.840 1.755 2.390 1.985 ;
        RECT  0.440 1.755 0.840 2.175 ;
        RECT  0.215 1.755 0.440 2.075 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 2.260 1.840 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 -0.400 3.300 0.400 ;
        RECT  2.780 -0.400 3.120 1.020 ;
        RECT  1.680 -0.400 2.780 0.400 ;
        RECT  1.340 -0.400 1.680 1.490 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 4.640 3.300 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  0.520 4.640 2.780 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR2X2

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2XL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.620 1.240 1.850 3.250 ;
        RECT  1.160 1.240 1.620 1.470 ;
        RECT  1.460 2.630 1.620 3.250 ;
        RECT  0.820 1.130 1.160 1.470 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.380 0.840 2.700 ;
        RECT  0.200 2.300 0.540 2.700 ;
        RECT  0.140 2.380 0.200 2.700 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.710 1.390 2.110 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 -0.400 1.980 0.400 ;
        RECT  1.460 -0.400 1.800 0.575 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 1.980 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NOR2X1

MACRO NAND4BBXL
    CLASS CORE ;
    FOREIGN NAND4BBXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 0.845 5.100 3.920 ;
        RECT  4.760 0.845 4.870 1.285 ;
        RECT  4.835 2.405 4.870 2.635 ;
        RECT  3.320 3.690 4.870 3.920 ;
        RECT  3.715 0.845 4.760 1.075 ;
        RECT  3.375 0.845 3.715 1.185 ;
        RECT  3.090 3.095 3.320 3.920 ;
        RECT  2.980 3.095 3.090 3.435 ;
        RECT  1.910 3.205 2.980 3.435 ;
        RECT  1.570 3.095 1.910 3.435 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.845 1.765 2.075 ;
        RECT  1.325 1.845 1.555 2.520 ;
        RECT  1.235 2.180 1.325 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.315 1.845 2.425 2.075 ;
        RECT  2.085 1.845 2.315 2.670 ;
        RECT  1.895 2.330 2.085 2.670 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.155 1.820 0.535 2.410 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.035 2.090 4.480 2.660 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 -0.400 5.280 0.400 ;
        RECT  4.760 -0.400 5.100 0.575 ;
        RECT  1.275 -0.400 4.760 0.400 ;
        RECT  0.455 -0.400 1.275 0.575 ;
        RECT  0.000 -0.400 0.455 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 4.640 5.280 5.440 ;
        RECT  3.610 4.465 4.060 5.440 ;
        RECT  2.615 4.640 3.610 5.440 ;
        RECT  2.275 4.465 2.615 5.440 ;
        RECT  1.315 4.640 2.275 5.440 ;
        RECT  0.865 4.465 1.315 5.440 ;
        RECT  0.000 4.640 0.865 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.410 3.095 4.640 3.435 ;
        RECT  4.080 1.305 4.420 1.840 ;
        RECT  3.790 3.095 4.410 3.325 ;
        RECT  3.790 1.610 4.080 1.840 ;
        RECT  3.560 1.610 3.790 3.325 ;
        RECT  3.355 1.760 3.560 2.100 ;
        RECT  2.785 1.340 3.015 2.670 ;
        RECT  0.995 1.340 2.785 1.570 ;
        RECT  2.675 2.330 2.785 2.670 ;
        RECT  0.765 1.340 0.995 3.335 ;
        RECT  0.520 1.340 0.765 1.570 ;
        RECT  0.520 3.105 0.765 3.335 ;
        RECT  0.180 1.230 0.520 1.570 ;
        RECT  0.180 3.105 0.520 3.445 ;
    END
END NAND4BBXL

MACRO NAND4BBX4
    CLASS CORE ;
    FOREIGN NAND4BBX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BBXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 1.820 12.400 3.220 ;
        RECT  12.060 0.805 12.360 3.955 ;
        RECT  12.020 0.805 12.060 1.290 ;
        RECT  12.020 1.820 12.060 3.220 ;
        RECT  8.515 3.655 12.060 3.955 ;
        RECT  8.800 0.805 12.020 1.105 ;
        RECT  8.600 0.630 8.800 1.105 ;
        RECT  8.260 0.630 8.600 1.440 ;
        RECT  1.735 3.655 8.515 3.935 ;
        RECT  3.720 0.870 8.260 1.150 ;
        RECT  3.380 0.630 3.720 1.440 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.530 2.180 10.640 2.520 ;
        RECT  10.300 2.180 10.530 3.425 ;
        RECT  6.160 3.195 10.300 3.425 ;
        RECT  5.820 3.085 6.160 3.425 ;
        RECT  1.765 3.195 5.820 3.425 ;
        RECT  1.680 2.965 1.765 3.425 ;
        RECT  1.535 2.180 1.680 3.425 ;
        RECT  1.450 2.180 1.535 3.195 ;
        RECT  1.340 2.180 1.450 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.905 2.180 9.960 2.520 ;
        RECT  9.620 2.180 9.905 2.660 ;
        RECT  9.610 2.405 9.620 2.660 ;
        RECT  9.455 2.405 9.610 2.965 ;
        RECT  9.380 2.430 9.455 2.965 ;
        RECT  7.115 2.735 9.380 2.965 ;
        RECT  6.775 2.625 7.115 2.965 ;
        RECT  5.200 2.625 6.775 2.855 ;
        RECT  4.860 2.625 5.200 2.965 ;
        RECT  2.425 2.735 4.860 2.965 ;
        RECT  2.195 2.180 2.425 2.965 ;
        RECT  2.020 2.180 2.195 2.520 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.360 2.010 11.740 2.700 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.155 1.820 0.535 2.410 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 -0.400 12.540 0.400 ;
        RECT  12.020 -0.400 12.360 0.575 ;
        RECT  11.040 -0.400 12.020 0.400 ;
        RECT  10.700 -0.400 11.040 0.575 ;
        RECT  6.160 -0.400 10.700 0.400 ;
        RECT  5.820 -0.400 6.160 0.575 ;
        RECT  1.280 -0.400 5.820 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.955 4.640 12.540 5.440 ;
        RECT  10.615 4.465 10.955 5.440 ;
        RECT  9.535 4.640 10.615 5.440 ;
        RECT  9.195 4.465 9.535 5.440 ;
        RECT  8.165 4.640 9.195 5.440 ;
        RECT  7.715 4.465 8.165 5.440 ;
        RECT  4.265 4.640 7.715 5.440 ;
        RECT  3.815 4.465 4.265 5.440 ;
        RECT  2.785 4.640 3.815 5.440 ;
        RECT  2.445 4.465 2.785 5.440 ;
        RECT  1.365 4.640 2.445 5.440 ;
        RECT  1.025 4.465 1.365 5.440 ;
        RECT  0.000 4.640 1.025 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.435 3.070 11.775 3.410 ;
        RECT  11.420 1.335 11.760 1.675 ;
        RECT  11.110 3.070 11.435 3.300 ;
        RECT  11.110 1.445 11.420 1.675 ;
        RECT  10.880 1.445 11.110 3.300 ;
        RECT  10.875 1.445 10.880 1.935 ;
        RECT  9.150 1.705 10.875 1.935 ;
        RECT  8.920 1.705 9.150 2.505 ;
        RECT  8.775 2.165 8.920 2.505 ;
        RECT  7.810 2.275 8.775 2.505 ;
        RECT  8.095 1.680 8.470 2.045 ;
        RECT  3.750 1.680 8.095 1.910 ;
        RECT  7.435 2.140 7.810 2.505 ;
        RECT  4.535 2.140 7.435 2.370 ;
        RECT  4.160 2.140 4.535 2.505 ;
        RECT  3.060 2.275 4.160 2.505 ;
        RECT  3.375 1.680 3.750 2.045 ;
        RECT  1.010 1.680 3.375 1.910 ;
        RECT  2.685 2.165 3.060 2.505 ;
        RECT  0.780 1.270 1.010 3.595 ;
        RECT  0.520 1.270 0.780 1.500 ;
        RECT  0.520 3.365 0.780 3.595 ;
        RECT  0.180 1.160 0.520 1.500 ;
        RECT  0.180 3.365 0.520 3.705 ;
    END
END NAND4BBX4

MACRO NAND4BBX2
    CLASS CORE ;
    FOREIGN NAND4BBX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BBXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.840 0.820 7.120 4.085 ;
        RECT  3.595 0.820 6.840 1.100 ;
        RECT  6.820 2.405 6.840 4.085 ;
        RECT  6.780 2.405 6.820 2.705 ;
        RECT  6.740 3.750 6.820 4.085 ;
        RECT  3.830 3.785 6.740 4.085 ;
        RECT  3.530 3.655 3.830 4.085 ;
        RECT  3.255 0.630 3.595 1.440 ;
        RECT  1.610 3.655 3.530 3.955 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.975 3.195 5.315 3.535 ;
        RECT  1.765 3.195 4.975 3.425 ;
        RECT  1.555 2.965 1.765 3.425 ;
        RECT  1.325 2.180 1.555 3.425 ;
        RECT  1.235 2.180 1.325 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.010 2.405 5.065 2.635 ;
        RECT  4.900 2.180 5.010 2.635 ;
        RECT  4.670 2.180 4.900 2.965 ;
        RECT  2.300 2.735 4.670 2.965 ;
        RECT  2.070 2.180 2.300 2.965 ;
        RECT  1.895 2.180 2.070 2.520 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.015 2.090 6.460 2.660 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.155 1.820 0.535 2.410 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.035 -0.400 7.260 0.400 ;
        RECT  5.695 -0.400 6.035 0.575 ;
        RECT  1.155 -0.400 5.695 0.400 ;
        RECT  0.335 -0.400 1.155 0.575 ;
        RECT  0.000 -0.400 0.335 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.830 4.640 7.260 5.440 ;
        RECT  6.305 4.465 6.830 5.440 ;
        RECT  4.140 4.640 6.305 5.440 ;
        RECT  3.690 4.465 4.140 5.440 ;
        RECT  2.660 4.640 3.690 5.440 ;
        RECT  2.320 4.465 2.660 5.440 ;
        RECT  1.240 4.640 2.320 5.440 ;
        RECT  0.900 4.465 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.380 1.330 6.610 1.670 ;
        RECT  5.775 1.385 6.380 1.670 ;
        RECT  5.775 3.195 5.885 3.535 ;
        RECT  5.545 1.385 5.775 3.535 ;
        RECT  4.355 1.685 5.545 1.915 ;
        RECT  4.125 1.685 4.355 2.505 ;
        RECT  3.980 2.160 4.125 2.505 ;
        RECT  2.935 2.275 3.980 2.505 ;
        RECT  3.250 1.680 3.625 2.045 ;
        RECT  0.995 1.680 3.250 1.910 ;
        RECT  2.560 2.165 2.935 2.505 ;
        RECT  0.765 1.270 0.995 3.065 ;
        RECT  0.520 1.270 0.765 1.500 ;
        RECT  0.520 2.835 0.765 3.065 ;
        RECT  0.180 1.160 0.520 1.500 ;
        RECT  0.180 2.835 0.520 3.645 ;
    END
END NAND4BBX2

MACRO NAND4BBX1
    CLASS CORE ;
    FOREIGN NAND4BBX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BBXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.065 2.405 5.155 3.920 ;
        RECT  4.925 0.845 5.065 3.920 ;
        RECT  4.835 0.845 4.925 2.635 ;
        RECT  3.310 3.690 4.925 3.920 ;
        RECT  4.760 0.845 4.835 1.285 ;
        RECT  3.635 0.845 4.760 1.075 ;
        RECT  3.295 0.845 3.635 1.185 ;
        RECT  3.080 3.115 3.310 3.920 ;
        RECT  2.970 3.115 3.080 3.525 ;
        RECT  2.780 3.170 2.970 3.525 ;
        RECT  2.195 3.170 2.780 3.400 ;
        RECT  1.950 3.115 2.195 3.400 ;
        RECT  1.610 3.115 1.950 3.455 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.845 1.765 2.075 ;
        RECT  1.325 1.845 1.555 2.520 ;
        RECT  1.235 2.180 1.325 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.300 1.845 2.425 2.075 ;
        RECT  2.070 1.845 2.300 2.670 ;
        RECT  1.895 2.330 2.070 2.670 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.155 1.820 0.535 2.410 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 2.090 4.530 2.430 ;
        RECT  4.035 2.090 4.480 2.660 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 -0.400 5.280 0.400 ;
        RECT  4.760 -0.400 5.100 0.575 ;
        RECT  1.190 -0.400 4.760 0.400 ;
        RECT  0.370 -0.400 1.190 0.575 ;
        RECT  0.000 -0.400 0.370 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 4.640 5.280 5.440 ;
        RECT  3.610 4.465 4.060 5.440 ;
        RECT  2.630 4.640 3.610 5.440 ;
        RECT  2.290 4.465 2.630 5.440 ;
        RECT  1.270 4.640 2.290 5.440 ;
        RECT  1.215 4.465 1.270 5.440 ;
        RECT  0.985 4.410 1.215 5.440 ;
        RECT  0.930 4.465 0.985 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.790 3.170 4.695 3.400 ;
        RECT  3.995 1.305 4.335 1.645 ;
        RECT  3.790 1.415 3.995 1.645 ;
        RECT  3.560 1.415 3.790 3.400 ;
        RECT  3.355 1.760 3.560 2.100 ;
        RECT  2.785 1.270 3.015 2.670 ;
        RECT  0.995 1.270 2.785 1.500 ;
        RECT  2.675 2.330 2.785 2.670 ;
        RECT  0.765 1.270 0.995 3.365 ;
        RECT  0.520 1.270 0.765 1.500 ;
        RECT  0.520 3.135 0.765 3.365 ;
        RECT  0.180 1.230 0.520 1.570 ;
        RECT  0.180 3.135 0.520 3.475 ;
    END
END NAND4BBX1

MACRO NAND4BXL
    CLASS CORE ;
    FOREIGN NAND4BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 3.525 3.085 3.755 ;
        RECT  2.420 1.060 2.760 1.400 ;
        RECT  2.300 1.170 2.420 1.400 ;
        RECT  2.300 3.525 2.405 3.945 ;
        RECT  2.070 1.170 2.300 3.945 ;
        RECT  1.765 3.605 2.070 3.945 ;
        RECT  1.080 3.715 1.765 3.945 ;
        RECT  0.740 3.605 1.080 3.945 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.280 1.845 0.600 2.520 ;
        RECT  0.215 1.845 0.280 2.515 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.775 1.380 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 1.820 1.840 2.235 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.145 2.295 3.820 2.740 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 -0.400 3.960 0.400 ;
        RECT  3.105 -0.400 3.445 0.575 ;
        RECT  0.520 -0.400 3.105 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.175 4.640 3.960 5.440 ;
        RECT  2.835 4.465 3.175 5.440 ;
        RECT  1.840 4.640 2.835 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.520 4.640 1.500 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.625 3.385 3.735 3.725 ;
        RECT  3.395 3.040 3.625 3.725 ;
        RECT  3.455 1.345 3.565 1.685 ;
        RECT  3.225 1.345 3.455 2.025 ;
        RECT  2.770 3.040 3.395 3.270 ;
        RECT  2.770 1.795 3.225 2.025 ;
        RECT  2.540 1.795 2.770 3.270 ;
    END
END NAND4BXL

MACRO NAND4BX4
    CLASS CORE ;
    FOREIGN NAND4BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.075 2.380 11.080 3.780 ;
        RECT  11.040 1.210 11.075 3.780 ;
        RECT  10.845 1.210 11.040 3.955 ;
        RECT  8.600 1.210 10.845 1.440 ;
        RECT  10.700 2.380 10.845 3.955 ;
        RECT  8.515 3.655 10.700 3.955 ;
        RECT  8.260 0.630 8.600 1.440 ;
        RECT  1.735 3.655 8.515 3.935 ;
        RECT  3.720 0.870 8.260 1.150 ;
        RECT  3.380 0.630 3.720 1.440 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.450 1.790 10.615 2.130 ;
        RECT  10.280 1.790 10.450 3.425 ;
        RECT  10.220 1.845 10.280 3.425 ;
        RECT  6.160 3.195 10.220 3.425 ;
        RECT  5.820 3.085 6.160 3.425 ;
        RECT  1.765 3.195 5.820 3.425 ;
        RECT  1.680 2.965 1.765 3.425 ;
        RECT  1.535 2.180 1.680 3.425 ;
        RECT  1.450 2.180 1.535 3.195 ;
        RECT  1.340 2.180 1.450 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.905 2.180 9.960 2.520 ;
        RECT  9.620 2.180 9.905 2.660 ;
        RECT  9.610 2.405 9.620 2.660 ;
        RECT  9.455 2.405 9.610 2.965 ;
        RECT  9.380 2.430 9.455 2.965 ;
        RECT  7.115 2.735 9.380 2.965 ;
        RECT  6.775 2.625 7.115 2.965 ;
        RECT  5.200 2.625 6.775 2.855 ;
        RECT  4.860 2.625 5.200 2.965 ;
        RECT  2.425 2.735 4.860 2.965 ;
        RECT  2.195 2.180 2.425 2.965 ;
        RECT  2.020 2.180 2.195 2.520 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 2.165 9.150 2.505 ;
        RECT  8.720 1.820 9.100 2.505 ;
        RECT  7.810 2.275 8.720 2.505 ;
        RECT  7.435 2.140 7.810 2.505 ;
        RECT  4.535 2.140 7.435 2.370 ;
        RECT  4.160 2.140 4.535 2.505 ;
        RECT  3.060 2.275 4.160 2.505 ;
        RECT  2.685 2.165 3.060 2.505 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.155 1.820 0.535 2.410 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.040 -0.400 11.880 0.400 ;
        RECT  10.700 -0.400 11.040 0.575 ;
        RECT  6.160 -0.400 10.700 0.400 ;
        RECT  5.820 -0.400 6.160 0.575 ;
        RECT  1.280 -0.400 5.820 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.955 4.640 11.880 5.440 ;
        RECT  10.615 4.465 10.955 5.440 ;
        RECT  9.535 4.640 10.615 5.440 ;
        RECT  9.195 4.465 9.535 5.440 ;
        RECT  8.165 4.640 9.195 5.440 ;
        RECT  7.715 4.465 8.165 5.440 ;
        RECT  4.265 4.640 7.715 5.440 ;
        RECT  3.815 4.465 4.265 5.440 ;
        RECT  2.785 4.640 3.815 5.440 ;
        RECT  2.445 4.465 2.785 5.440 ;
        RECT  1.365 4.640 2.445 5.440 ;
        RECT  1.025 4.465 1.365 5.440 ;
        RECT  0.000 4.640 1.025 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.095 1.680 8.470 2.045 ;
        RECT  3.750 1.680 8.095 1.910 ;
        RECT  3.375 1.680 3.750 2.045 ;
        RECT  1.010 1.680 3.375 1.910 ;
        RECT  0.780 1.270 1.010 3.595 ;
        RECT  0.520 1.270 0.780 1.500 ;
        RECT  0.520 3.365 0.780 3.595 ;
        RECT  0.180 1.160 0.520 1.500 ;
        RECT  0.180 3.365 0.520 3.705 ;
    END
END NAND4BX4

MACRO NAND4BX2
    CLASS CORE ;
    FOREIGN NAND4BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.380 0.820 6.385 2.660 ;
        RECT  6.105 0.820 6.380 4.085 ;
        RECT  6.080 0.820 6.105 1.285 ;
        RECT  6.080 2.370 6.105 4.085 ;
        RECT  3.620 0.820 6.080 1.100 ;
        RECT  3.830 3.785 6.080 4.085 ;
        RECT  3.530 3.655 3.830 4.085 ;
        RECT  3.280 0.630 3.620 1.440 ;
        RECT  1.610 3.655 3.530 3.955 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.975 3.195 5.315 3.535 ;
        RECT  1.765 3.195 4.975 3.425 ;
        RECT  1.555 2.965 1.765 3.425 ;
        RECT  1.535 2.180 1.555 3.425 ;
        RECT  1.325 2.180 1.535 3.195 ;
        RECT  1.245 2.180 1.325 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.050 2.405 5.065 2.635 ;
        RECT  4.940 2.180 5.050 2.635 ;
        RECT  4.710 2.180 4.940 2.965 ;
        RECT  2.300 2.735 4.710 2.965 ;
        RECT  2.070 2.180 2.300 2.965 ;
        RECT  1.910 2.180 2.070 2.520 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.355 1.845 4.405 2.075 ;
        RECT  4.100 1.820 4.355 2.505 ;
        RECT  3.980 2.160 4.100 2.505 ;
        RECT  2.935 2.275 3.980 2.505 ;
        RECT  2.560 2.165 2.935 2.505 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.155 1.820 0.535 2.410 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.060 -0.400 6.600 0.400 ;
        RECT  5.720 -0.400 6.060 0.575 ;
        RECT  1.180 -0.400 5.720 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 4.640 6.600 5.440 ;
        RECT  3.690 4.465 4.140 5.440 ;
        RECT  2.660 4.640 3.690 5.440 ;
        RECT  2.320 4.465 2.660 5.440 ;
        RECT  1.240 4.640 2.320 5.440 ;
        RECT  1.185 4.465 1.240 5.440 ;
        RECT  0.955 4.410 1.185 5.440 ;
        RECT  0.900 4.465 0.955 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.250 1.680 3.625 2.045 ;
        RECT  1.005 1.680 3.250 1.910 ;
        RECT  0.775 1.270 1.005 3.355 ;
        RECT  0.520 1.270 0.775 1.500 ;
        RECT  0.520 3.125 0.775 3.355 ;
        RECT  0.180 1.160 0.520 1.500 ;
        RECT  0.180 3.070 0.520 3.410 ;
    END
END NAND4BX2

MACRO NAND4BX1
    CLASS CORE ;
    FOREIGN NAND4BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 2.405 4.495 3.920 ;
        RECT  4.265 0.845 4.405 3.920 ;
        RECT  4.175 0.845 4.265 2.635 ;
        RECT  2.650 3.690 4.265 3.920 ;
        RECT  4.100 0.845 4.175 1.285 ;
        RECT  2.975 0.845 4.100 1.075 ;
        RECT  2.635 0.845 2.975 1.185 ;
        RECT  2.420 3.095 2.650 3.920 ;
        RECT  2.310 3.095 2.420 3.525 ;
        RECT  2.120 3.205 2.310 3.525 ;
        RECT  1.290 3.205 2.120 3.435 ;
        RECT  0.950 3.095 1.290 3.435 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 1.845 1.105 2.075 ;
        RECT  0.665 1.845 0.895 2.520 ;
        RECT  0.575 2.065 0.665 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 1.845 1.765 2.075 ;
        RECT  1.575 1.845 1.655 2.615 ;
        RECT  1.425 1.845 1.575 2.670 ;
        RECT  1.235 2.330 1.425 2.670 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 2.330 2.640 2.795 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 2.090 3.870 2.430 ;
        RECT  3.375 2.090 3.820 2.660 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 -0.400 4.620 0.400 ;
        RECT  4.100 -0.400 4.440 0.575 ;
        RECT  0.535 -0.400 4.100 0.400 ;
        RECT  0.195 -0.400 0.535 0.575 ;
        RECT  0.000 -0.400 0.195 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 4.640 4.620 5.440 ;
        RECT  2.950 4.465 3.400 5.440 ;
        RECT  1.970 4.640 2.950 5.440 ;
        RECT  1.630 4.465 1.970 5.440 ;
        RECT  0.620 4.640 1.630 5.440 ;
        RECT  0.280 4.465 0.620 5.440 ;
        RECT  0.000 4.640 0.280 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.695 3.095 4.035 3.435 ;
        RECT  3.130 3.095 3.695 3.325 ;
        RECT  3.525 1.305 3.675 1.645 ;
        RECT  3.335 1.305 3.525 1.700 ;
        RECT  3.295 1.360 3.335 1.700 ;
        RECT  3.130 1.470 3.295 1.700 ;
        RECT  2.900 1.470 3.130 3.325 ;
        RECT  2.695 1.760 2.900 2.100 ;
    END
END NAND4BX1

MACRO NAND4XL
    CLASS CORE ;
    FOREIGN NAND4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.420 1.245 2.975 1.585 ;
        RECT  2.170 3.095 2.510 3.435 ;
        RECT  1.765 1.355 2.420 1.585 ;
        RECT  1.765 3.095 2.170 3.325 ;
        RECT  1.535 1.355 1.765 3.325 ;
        RECT  1.130 3.095 1.535 3.325 ;
        RECT  0.790 3.095 1.130 3.435 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.345 0.645 2.685 ;
        RECT  0.290 1.845 0.520 2.685 ;
        RECT  0.215 1.845 0.290 2.075 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 2.345 1.270 2.685 ;
        RECT  0.980 1.845 1.210 2.685 ;
        RECT  0.875 1.845 0.980 2.075 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.285 1.845 2.425 2.075 ;
        RECT  2.055 1.845 2.285 2.685 ;
        RECT  1.995 2.345 2.055 2.685 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 1.845 3.085 2.075 ;
        RECT  2.780 1.845 3.070 2.685 ;
        RECT  2.730 2.345 2.780 2.685 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 -0.400 3.300 0.400 ;
        RECT  0.195 -0.400 0.535 0.575 ;
        RECT  0.000 -0.400 0.195 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 4.640 3.300 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  2.085 4.640 2.780 5.440 ;
        RECT  1.730 4.465 2.085 5.440 ;
        RECT  0.520 4.640 1.730 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NAND4XL

MACRO NAND4X4
    CLASS CORE ;
    FOREIGN NAND4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4XL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.420 0.805 10.485 2.685 ;
        RECT  10.380 0.805 10.420 3.780 ;
        RECT  10.185 0.805 10.380 3.955 ;
        RECT  10.040 0.805 10.185 1.290 ;
        RECT  10.040 2.380 10.185 3.955 ;
        RECT  8.140 0.805 10.040 1.105 ;
        RECT  7.855 3.655 10.040 3.955 ;
        RECT  7.940 0.630 8.140 1.105 ;
        RECT  7.600 0.630 7.940 1.440 ;
        RECT  1.075 3.655 7.855 3.935 ;
        RECT  3.060 0.870 7.600 1.150 ;
        RECT  2.720 0.630 3.060 1.440 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.790 1.790 9.955 2.130 ;
        RECT  9.620 1.790 9.790 3.425 ;
        RECT  9.560 1.845 9.620 3.425 ;
        RECT  5.500 3.195 9.560 3.425 ;
        RECT  5.160 3.085 5.500 3.425 ;
        RECT  1.105 3.195 5.160 3.425 ;
        RECT  1.020 2.965 1.105 3.425 ;
        RECT  0.875 2.180 1.020 3.425 ;
        RECT  0.790 2.180 0.875 3.195 ;
        RECT  0.680 2.180 0.790 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.245 2.180 9.300 2.520 ;
        RECT  8.960 2.180 9.245 2.660 ;
        RECT  8.950 2.405 8.960 2.660 ;
        RECT  8.795 2.405 8.950 2.965 ;
        RECT  8.720 2.430 8.795 2.965 ;
        RECT  6.455 2.735 8.720 2.965 ;
        RECT  6.115 2.625 6.455 2.965 ;
        RECT  4.540 2.625 6.115 2.855 ;
        RECT  4.200 2.625 4.540 2.965 ;
        RECT  1.765 2.735 4.200 2.965 ;
        RECT  1.535 2.180 1.765 2.965 ;
        RECT  1.360 2.180 1.535 2.520 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.440 2.165 8.490 2.505 ;
        RECT  8.060 1.820 8.440 2.505 ;
        RECT  7.150 2.275 8.060 2.505 ;
        RECT  6.775 2.140 7.150 2.505 ;
        RECT  3.875 2.140 6.775 2.370 ;
        RECT  3.500 2.140 3.875 2.505 ;
        RECT  2.400 2.275 3.500 2.505 ;
        RECT  2.025 2.165 2.400 2.505 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.435 1.680 7.810 2.045 ;
        RECT  3.090 1.680 7.435 1.910 ;
        RECT  2.715 1.680 3.090 2.045 ;
        RECT  1.840 1.680 2.715 1.910 ;
        RECT  1.610 1.285 1.840 1.910 ;
        RECT  1.535 1.285 1.610 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.380 -0.400 11.220 0.400 ;
        RECT  10.040 -0.400 10.380 0.575 ;
        RECT  5.500 -0.400 10.040 0.400 ;
        RECT  5.160 -0.400 5.500 0.575 ;
        RECT  0.620 -0.400 5.160 0.400 ;
        RECT  0.280 -0.400 0.620 0.575 ;
        RECT  0.000 -0.400 0.280 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.295 4.640 11.220 5.440 ;
        RECT  9.955 4.465 10.295 5.440 ;
        RECT  8.875 4.640 9.955 5.440 ;
        RECT  8.535 4.465 8.875 5.440 ;
        RECT  7.505 4.640 8.535 5.440 ;
        RECT  7.055 4.465 7.505 5.440 ;
        RECT  3.605 4.640 7.055 5.440 ;
        RECT  3.155 4.465 3.605 5.440 ;
        RECT  2.125 4.640 3.155 5.440 ;
        RECT  1.785 4.465 2.125 5.440 ;
        RECT  0.705 4.640 1.785 5.440 ;
        RECT  0.365 4.465 0.705 5.440 ;
        RECT  0.000 4.640 0.365 5.440 ;
        END
    END VDD
END NAND4X4

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 0.820 5.725 2.660 ;
        RECT  5.445 0.820 5.720 4.085 ;
        RECT  5.420 0.820 5.445 1.285 ;
        RECT  5.420 2.370 5.445 4.085 ;
        RECT  2.960 0.820 5.420 1.100 ;
        RECT  3.170 3.785 5.420 4.085 ;
        RECT  2.870 3.655 3.170 4.085 ;
        RECT  2.620 0.630 2.960 1.440 ;
        RECT  0.950 3.655 2.870 3.955 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.315 3.195 4.655 3.535 ;
        RECT  1.105 3.195 4.315 3.425 ;
        RECT  0.895 2.965 1.105 3.425 ;
        RECT  0.875 2.180 0.895 3.425 ;
        RECT  0.665 2.180 0.875 3.195 ;
        RECT  0.555 2.180 0.665 2.520 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 2.180 4.430 2.520 ;
        RECT  4.320 2.180 4.405 2.635 ;
        RECT  4.090 2.180 4.320 2.965 ;
        RECT  1.640 2.735 4.090 2.965 ;
        RECT  1.410 2.180 1.640 2.965 ;
        RECT  1.235 2.180 1.410 2.520 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 1.845 3.775 2.505 ;
        RECT  2.275 2.275 3.400 2.505 ;
        RECT  1.900 2.165 2.275 2.505 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.590 1.685 2.965 2.045 ;
        RECT  1.840 1.685 2.590 1.915 ;
        RECT  1.610 1.285 1.840 1.915 ;
        RECT  1.535 1.285 1.610 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.400 -0.400 5.940 0.400 ;
        RECT  5.060 -0.400 5.400 0.575 ;
        RECT  0.520 -0.400 5.060 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.480 4.640 5.940 5.440 ;
        RECT  3.030 4.465 3.480 5.440 ;
        RECT  2.000 4.640 3.030 5.440 ;
        RECT  1.660 4.465 2.000 5.440 ;
        RECT  0.580 4.640 1.660 5.440 ;
        RECT  0.240 4.465 0.580 5.440 ;
        RECT  0.000 4.640 0.240 5.440 ;
        END
    END VDD
END NAND4X2

MACRO NAND4X1
    CLASS CORE ;
    FOREIGN NAND4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.995 1.295 3.170 3.325 ;
        RECT  2.940 0.715 2.995 3.325 ;
        RECT  2.655 0.715 2.940 1.525 ;
        RECT  2.780 2.965 2.940 3.325 ;
        RECT  2.500 3.095 2.780 3.325 ;
        RECT  2.160 3.095 2.500 3.435 ;
        RECT  1.140 3.095 2.160 3.325 ;
        RECT  0.800 3.095 1.140 3.435 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.330 0.770 2.670 ;
        RECT  0.290 1.845 0.520 2.670 ;
        RECT  0.215 1.845 0.290 2.075 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 2.330 1.485 2.670 ;
        RECT  1.000 1.845 1.230 2.670 ;
        RECT  0.875 1.845 1.000 2.075 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.910 2.405 2.500 2.780 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 1.760 2.705 2.100 ;
        RECT  1.535 1.845 2.365 2.075 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 -0.400 3.300 0.400 ;
        RECT  0.195 -0.400 0.535 1.100 ;
        RECT  0.000 -0.400 0.195 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 4.640 3.300 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  2.080 4.640 2.780 5.440 ;
        RECT  1.740 4.465 2.080 5.440 ;
        RECT  0.520 4.640 1.740 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NAND4X1

MACRO NAND3BXL
    CLASS CORE ;
    FOREIGN NAND3BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 0.665 3.160 4.375 ;
        RECT  2.720 0.665 2.930 0.895 ;
        RECT  2.855 2.940 2.930 4.375 ;
        RECT  2.780 2.940 2.855 3.585 ;
        RECT  2.760 4.145 2.855 4.375 ;
        RECT  1.840 3.355 2.780 3.585 ;
        RECT  1.500 3.300 1.840 3.640 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 2.550 1.440 3.020 ;
        RECT  1.210 2.550 1.215 3.220 ;
        RECT  0.800 2.790 1.210 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.590 2.130 2.100 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.540 0.520 2.100 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 -0.400 3.300 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 4.640 3.300 5.440 ;
        RECT  2.060 4.465 2.400 5.440 ;
        RECT  1.180 4.640 2.060 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.465 1.125 2.695 2.550 ;
        RECT  0.980 1.125 2.465 1.355 ;
        RECT  0.750 1.080 0.980 2.560 ;
        RECT  0.180 1.080 0.750 1.310 ;
        RECT  0.465 2.330 0.750 2.560 ;
        RECT  0.465 3.210 0.520 3.550 ;
        RECT  0.235 2.330 0.465 3.550 ;
        RECT  0.180 3.210 0.235 3.550 ;
    END
END NAND3BXL

MACRO NAND3BX4
    CLASS CORE ;
    FOREIGN NAND3BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3BXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.850 0.835 7.080 3.170 ;
        RECT  6.700 0.835 6.850 1.290 ;
        RECT  6.460 2.940 6.850 3.170 ;
        RECT  3.200 0.835 6.700 1.065 ;
        RECT  6.255 2.940 6.460 4.340 ;
        RECT  6.080 2.890 6.255 4.340 ;
        RECT  5.725 2.890 6.080 3.400 ;
        RECT  3.545 3.170 5.725 3.400 ;
        RECT  3.205 3.115 3.545 3.455 ;
        RECT  3.085 3.115 3.205 3.400 ;
        RECT  2.860 0.700 3.200 1.065 ;
        RECT  2.125 3.170 3.085 3.400 ;
        RECT  1.785 3.115 2.125 3.455 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 3.845 4.820 4.185 ;
        RECT  1.440 3.900 4.480 4.130 ;
        RECT  1.440 1.845 1.765 2.100 ;
        RECT  1.210 1.845 1.440 4.130 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.405 2.130 5.745 2.550 ;
        RECT  4.480 2.130 5.405 2.360 ;
        RECT  4.110 2.130 4.480 2.660 ;
        RECT  3.770 2.075 4.110 2.660 ;
        RECT  3.745 2.380 3.770 2.660 ;
        RECT  2.400 2.430 3.745 2.660 ;
        RECT  2.060 2.425 2.400 2.765 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.170 1.725 0.510 2.365 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 -0.400 7.260 0.400 ;
        RECT  4.760 -0.400 5.100 0.575 ;
        RECT  1.300 -0.400 4.760 0.400 ;
        RECT  0.960 -0.400 1.300 0.575 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.920 4.640 7.260 5.440 ;
        RECT  6.690 3.740 6.920 5.440 ;
        RECT  5.545 4.640 6.690 5.440 ;
        RECT  5.205 3.740 5.545 5.440 ;
        RECT  4.225 4.640 5.205 5.440 ;
        RECT  3.885 4.465 4.225 5.440 ;
        RECT  2.835 4.640 3.885 5.440 ;
        RECT  2.495 4.465 2.835 5.440 ;
        RECT  1.315 4.640 2.495 5.440 ;
        RECT  0.975 4.465 1.315 5.440 ;
        RECT  0.000 4.640 0.975 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.445 1.850 6.615 2.330 ;
        RECT  6.385 1.325 6.445 2.330 ;
        RECT  6.215 1.325 6.385 2.080 ;
        RECT  3.080 1.325 6.215 1.555 ;
        RECT  2.740 1.325 3.080 2.085 ;
        RECT  0.980 1.325 2.740 1.555 ;
        RECT  0.750 1.050 0.980 3.130 ;
        RECT  0.520 1.050 0.750 1.280 ;
        RECT  0.520 2.900 0.750 3.130 ;
        RECT  0.180 0.940 0.520 1.280 ;
        RECT  0.180 2.900 0.520 3.240 ;
    END
END NAND3BX4

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.455 2.895 2.795 3.235 ;
        RECT  2.140 0.690 2.480 1.030 ;
        RECT  2.425 2.895 2.455 3.220 ;
        RECT  1.535 2.940 2.425 3.220 ;
        RECT  1.110 0.745 2.140 0.975 ;
        RECT  1.405 2.895 1.535 3.220 ;
        RECT  1.110 2.895 1.405 3.235 ;
        RECT  1.065 0.745 1.110 3.235 ;
        RECT  0.880 0.745 1.065 3.220 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 1.940 3.950 2.280 ;
        RECT  3.665 1.940 3.895 3.700 ;
        RECT  3.610 1.940 3.665 2.280 ;
        RECT  0.650 3.470 3.665 3.700 ;
        RECT  0.420 1.845 0.650 3.700 ;
        RECT  0.310 1.845 0.420 2.405 ;
        RECT  0.215 1.845 0.310 2.075 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 2.130 3.280 2.470 ;
        RECT  2.780 1.820 3.160 2.535 ;
        RECT  1.680 2.305 2.780 2.535 ;
        RECT  1.340 2.160 1.680 2.535 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.120 1.960 5.140 2.495 ;
        RECT  4.780 1.820 5.120 2.495 ;
        RECT  4.760 1.960 4.780 2.495 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 -0.400 5.280 0.400 ;
        RECT  4.320 -0.400 4.380 0.575 ;
        RECT  3.980 -0.400 4.320 1.100 ;
        RECT  0.580 -0.400 3.980 0.400 ;
        RECT  0.240 -0.400 0.580 1.100 ;
        RECT  0.000 -0.400 0.240 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 4.640 5.280 5.440 ;
        RECT  3.990 3.935 4.330 5.440 ;
        RECT  2.115 4.640 3.990 5.440 ;
        RECT  1.775 3.935 2.115 5.440 ;
        RECT  0.725 4.640 1.775 5.440 ;
        RECT  0.385 3.935 0.725 5.440 ;
        RECT  0.000 4.640 0.385 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.760 1.170 5.100 1.590 ;
        RECT  4.760 2.950 5.100 3.290 ;
        RECT  4.530 1.360 4.760 1.590 ;
        RECT  4.530 2.950 4.760 3.180 ;
        RECT  4.300 1.360 4.530 3.180 ;
        RECT  2.480 1.360 4.300 1.590 ;
        RECT  2.250 1.360 2.480 2.060 ;
        RECT  2.140 1.720 2.250 2.060 ;
    END
END NAND3BX2

MACRO NAND3BX1
    CLASS CORE ;
    FOREIGN NAND3BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3BXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 0.665 3.160 4.375 ;
        RECT  2.720 0.665 2.930 0.895 ;
        RECT  2.855 3.500 2.930 4.375 ;
        RECT  1.840 3.500 2.855 3.730 ;
        RECT  2.760 4.145 2.855 4.375 ;
        RECT  1.500 3.500 1.840 3.840 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 2.490 1.440 3.195 ;
        RECT  0.875 2.795 1.210 3.195 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.740 2.080 2.100 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.540 0.520 2.100 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 3.300 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 4.640 3.300 5.440 ;
        RECT  2.060 4.465 2.400 5.440 ;
        RECT  1.180 4.640 2.060 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.465 1.125 2.695 2.540 ;
        RECT  0.980 1.125 2.465 1.355 ;
        RECT  0.750 1.080 0.980 2.560 ;
        RECT  0.180 1.080 0.750 1.310 ;
        RECT  0.465 2.330 0.750 2.560 ;
        RECT  0.465 3.585 0.520 3.925 ;
        RECT  0.235 2.330 0.465 3.925 ;
        RECT  0.180 3.585 0.235 3.925 ;
    END
END NAND3BX1

MACRO NAND3XL
    CLASS CORE ;
    FOREIGN NAND3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 1.055 2.460 3.285 ;
        RECT  2.120 1.055 2.230 1.395 ;
        RECT  2.120 2.860 2.230 3.285 ;
        RECT  1.050 3.055 2.120 3.285 ;
        RECT  0.710 3.000 1.050 3.340 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.045 0.520 2.660 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.820 1.315 2.590 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 2.250 1.995 2.590 ;
        RECT  1.655 1.285 1.885 2.590 ;
        RECT  1.535 1.285 1.655 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.400 2.640 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.720 4.640 2.640 5.440 ;
        RECT  0.450 4.465 1.720 5.440 ;
        RECT  0.000 4.640 0.450 5.440 ;
        END
    END VDD
END NAND3XL

MACRO NAND3X4
    CLASS CORE ;
    FOREIGN NAND3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.260 0.665 6.280 1.475 ;
        RECT  6.030 0.665 6.260 3.125 ;
        RECT  5.940 0.665 6.030 1.475 ;
        RECT  5.535 2.895 6.030 3.125 ;
        RECT  5.720 0.665 5.940 1.040 ;
        RECT  2.480 0.810 5.720 1.040 ;
        RECT  5.195 2.895 5.535 3.235 ;
        RECT  1.160 2.895 2.825 3.235 ;
        RECT  1.180 0.700 2.480 1.040 ;
        RECT  1.160 0.700 1.180 2.100 ;
        RECT  0.820 0.700 1.160 3.235 ;
        RECT  0.800 0.700 0.820 2.100 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.025 2.215 4.080 2.555 ;
        RECT  3.795 2.215 4.025 3.695 ;
        RECT  3.740 2.215 3.795 2.555 ;
        RECT  0.570 3.465 3.795 3.695 ;
        RECT  0.340 1.845 0.570 3.695 ;
        RECT  0.215 1.845 0.340 2.405 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.005 2.075 5.115 2.480 ;
        RECT  4.775 1.755 5.005 2.480 ;
        RECT  3.400 1.755 4.775 1.985 ;
        RECT  3.060 1.750 3.400 2.090 ;
        RECT  3.010 1.755 3.060 2.090 ;
        RECT  2.780 1.755 3.010 2.525 ;
        RECT  1.750 2.295 2.780 2.525 ;
        RECT  1.410 2.160 1.750 2.525 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.670 1.790 5.790 2.480 ;
        RECT  5.450 1.270 5.670 2.480 ;
        RECT  5.440 1.270 5.450 2.095 ;
        RECT  2.480 1.270 5.440 1.500 ;
        RECT  2.250 1.270 2.480 2.065 ;
        RECT  2.140 1.725 2.250 2.065 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 -0.400 6.600 0.400 ;
        RECT  4.040 -0.400 4.380 0.575 ;
        RECT  0.570 -0.400 4.040 0.400 ;
        RECT  0.230 -0.400 0.570 1.100 ;
        RECT  0.000 -0.400 0.230 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.215 4.640 6.600 5.440 ;
        RECT  5.875 3.935 6.215 5.440 ;
        RECT  4.855 4.640 5.875 5.440 ;
        RECT  4.515 3.935 4.855 5.440 ;
        RECT  3.505 4.640 4.515 5.440 ;
        RECT  3.165 3.935 3.505 5.440 ;
        RECT  2.115 4.640 3.165 5.440 ;
        RECT  1.775 3.935 2.115 5.440 ;
        RECT  0.725 4.640 1.775 5.440 ;
        RECT  0.385 3.935 0.725 5.440 ;
        RECT  0.000 4.640 0.385 5.440 ;
        END
    END VDD
END NAND3X4

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.455 2.895 2.795 3.235 ;
        RECT  2.140 0.690 2.480 1.030 ;
        RECT  2.425 2.895 2.455 3.195 ;
        RECT  1.840 2.965 2.425 3.195 ;
        RECT  1.110 0.800 2.140 1.030 ;
        RECT  1.535 2.940 1.840 3.235 ;
        RECT  1.110 2.895 1.535 3.235 ;
        RECT  1.065 0.800 1.110 3.235 ;
        RECT  0.880 0.800 1.065 3.195 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 2.405 3.950 2.965 ;
        RECT  3.665 2.405 3.895 3.700 ;
        RECT  3.610 2.405 3.665 2.965 ;
        RECT  0.650 3.470 3.665 3.700 ;
        RECT  0.595 1.930 0.650 3.700 ;
        RECT  0.420 1.845 0.595 3.700 ;
        RECT  0.310 1.845 0.420 2.405 ;
        RECT  0.215 1.845 0.310 2.075 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.225 2.070 3.280 2.470 ;
        RECT  3.085 1.820 3.225 2.470 ;
        RECT  2.780 1.820 3.085 2.535 ;
        RECT  1.680 2.305 2.780 2.535 ;
        RECT  1.340 2.160 1.680 2.535 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.140 1.260 2.480 2.060 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 -0.400 4.620 0.400 ;
        RECT  4.040 -0.400 4.380 0.575 ;
        RECT  0.580 -0.400 4.040 0.400 ;
        RECT  0.240 -0.400 0.580 0.575 ;
        RECT  0.000 -0.400 0.240 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 4.640 4.620 5.440 ;
        RECT  1.775 3.935 2.115 5.440 ;
        RECT  0.725 4.640 1.775 5.440 ;
        RECT  0.385 3.935 0.725 5.440 ;
        RECT  0.000 4.640 0.385 5.440 ;
        END
    END VDD
END NAND3X2

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 2.920 2.470 3.410 ;
        RECT  2.230 0.700 2.460 3.410 ;
        RECT  2.120 0.700 2.230 1.290 ;
        RECT  2.190 2.920 2.230 3.410 ;
        RECT  2.120 3.070 2.190 3.410 ;
        RECT  1.105 3.125 2.120 3.355 ;
        RECT  0.765 3.070 1.105 3.410 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.190 1.785 0.530 2.480 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.285 1.315 2.840 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 2.105 1.995 2.445 ;
        RECT  1.655 1.285 1.885 2.445 ;
        RECT  1.535 1.285 1.655 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 -0.400 2.640 0.400 ;
        RECT  0.240 -0.400 0.580 0.575 ;
        RECT  0.000 -0.400 0.240 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 4.640 2.640 5.440 ;
        RECT  0.180 4.465 1.820 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NAND3X1

MACRO NAND2BXL
    CLASS CORE ;
    FOREIGN NAND2BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 1.285 2.495 3.550 ;
        RECT  2.265 1.030 2.440 3.550 ;
        RECT  2.100 1.030 2.265 1.515 ;
        RECT  1.840 3.320 2.265 3.550 ;
        RECT  1.535 1.285 2.100 1.515 ;
        RECT  1.500 3.265 1.840 3.605 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.420 1.930 1.475 2.285 ;
        RECT  0.875 1.845 1.420 2.285 ;
        RECT  0.800 1.930 0.875 2.285 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.210 3.785 0.740 4.340 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 4.640 2.640 5.440 ;
        RECT  1.420 4.465 2.400 5.440 ;
        RECT  0.000 4.640 1.420 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.795 2.575 2.025 3.035 ;
        RECT  0.520 2.805 1.795 3.035 ;
        RECT  0.465 1.150 0.520 1.490 ;
        RECT  0.465 2.805 0.520 3.450 ;
        RECT  0.235 1.150 0.465 3.450 ;
        RECT  0.180 1.150 0.235 1.490 ;
        RECT  0.180 3.110 0.235 3.450 ;
    END
END NAND2BXL

MACRO NAND2BX4
    CLASS CORE ;
    FOREIGN NAND2BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.120 1.030 5.140 2.660 ;
        RECT  4.780 1.030 5.120 3.350 ;
        RECT  4.760 1.030 4.780 2.660 ;
        RECT  1.495 3.010 4.780 3.350 ;
        RECT  2.540 1.375 4.760 1.675 ;
        RECT  2.200 1.190 2.540 1.675 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.385 3.715 2.780 ;
        RECT  1.810 2.550 3.085 2.780 ;
        RECT  1.600 2.405 1.810 2.780 ;
        RECT  1.260 2.385 1.600 2.780 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.170 2.020 0.510 2.660 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 -0.400 5.280 0.400 ;
        RECT  3.480 -0.400 3.820 1.130 ;
        RECT  1.280 -0.400 3.480 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.040 4.640 5.280 5.440 ;
        RECT  4.700 3.595 5.040 5.440 ;
        RECT  3.755 4.640 4.700 5.440 ;
        RECT  3.415 3.595 3.755 5.440 ;
        RECT  2.475 4.640 3.415 5.440 ;
        RECT  2.135 3.595 2.475 5.440 ;
        RECT  1.195 4.640 2.135 5.440 ;
        RECT  0.855 3.645 1.195 5.440 ;
        RECT  0.000 4.640 0.855 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.300 1.920 4.530 2.725 ;
        RECT  2.530 1.920 4.300 2.150 ;
        RECT  2.190 1.920 2.530 2.320 ;
        RECT  0.980 1.920 2.190 2.150 ;
        RECT  0.750 1.280 0.980 3.240 ;
        RECT  0.520 1.280 0.750 1.510 ;
        RECT  0.520 3.010 0.750 3.240 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  0.180 3.010 0.520 3.350 ;
    END
END NAND2BX4

MACRO NAND2BX2
    CLASS CORE ;
    FOREIGN NAND2BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.610 1.690 3.840 3.235 ;
        RECT  3.160 1.690 3.610 1.920 ;
        RECT  3.220 2.940 3.610 3.235 ;
        RECT  2.880 2.900 3.220 3.240 ;
        RECT  3.155 1.515 3.160 1.920 ;
        RECT  2.925 1.330 3.155 1.920 ;
        RECT  2.500 1.330 2.925 1.560 ;
        RECT  2.780 2.940 2.880 3.235 ;
        RECT  2.195 3.005 2.780 3.235 ;
        RECT  2.160 1.220 2.500 1.560 ;
        RECT  1.940 2.950 2.195 3.235 ;
        RECT  1.600 2.950 1.940 3.290 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 2.305 3.380 2.670 ;
        RECT  1.680 2.405 3.070 2.635 ;
        RECT  1.340 2.350 1.680 2.690 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.170 1.900 0.510 2.635 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 3.960 0.400 ;
        RECT  3.440 -0.400 3.780 1.230 ;
        RECT  1.180 -0.400 3.440 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 4.640 3.960 5.440 ;
        RECT  1.270 4.465 3.780 5.440 ;
        RECT  0.000 4.640 1.270 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.300 1.820 2.640 2.160 ;
        RECT  0.980 1.875 2.300 2.105 ;
        RECT  0.750 1.305 0.980 3.180 ;
        RECT  0.520 1.305 0.750 1.545 ;
        RECT  0.520 2.950 0.750 3.180 ;
        RECT  0.180 1.170 0.520 1.545 ;
        RECT  0.180 2.950 0.520 3.290 ;
        RECT  0.175 1.225 0.180 1.545 ;
    END
END NAND2BX2

MACRO NAND2BX1
    CLASS CORE ;
    FOREIGN NAND2BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2BXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 1.215 2.440 3.395 ;
        RECT  2.100 1.215 2.210 1.555 ;
        RECT  1.500 3.165 2.210 3.395 ;
        RECT  1.760 1.260 2.100 1.540 ;
        RECT  1.535 1.285 1.760 1.515 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.420 1.935 1.475 2.290 ;
        RECT  0.875 1.845 1.420 2.290 ;
        RECT  0.800 1.935 0.875 2.290 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.210 3.785 0.740 4.340 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 4.640 2.640 5.440 ;
        RECT  1.420 4.465 2.400 5.440 ;
        RECT  0.000 4.640 1.420 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.745 2.540 1.975 2.915 ;
        RECT  0.465 2.540 1.745 2.770 ;
        RECT  0.465 1.150 0.520 1.490 ;
        RECT  0.465 3.110 0.520 3.450 ;
        RECT  0.235 1.150 0.465 3.450 ;
        RECT  0.180 1.150 0.235 1.490 ;
        RECT  0.180 3.110 0.235 3.450 ;
    END
END NAND2BX1

MACRO NAND2XL
    CLASS CORE ;
    FOREIGN NAND2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 1.235 1.820 3.235 ;
        RECT  1.765 1.180 1.800 3.235 ;
        RECT  1.590 1.180 1.765 3.350 ;
        RECT  1.460 1.180 1.590 1.520 ;
        RECT  1.490 2.920 1.590 3.350 ;
        RECT  1.170 3.120 1.490 3.350 ;
        RECT  0.830 3.120 1.170 3.460 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.100 0.520 2.710 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 2.075 1.360 2.620 ;
        RECT  1.020 1.845 1.250 2.620 ;
        RECT  0.875 1.845 1.020 2.075 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.400 1.980 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.060 4.640 1.980 5.440 ;
        RECT  0.490 4.465 1.060 5.440 ;
        RECT  0.000 4.640 0.490 5.440 ;
        END
    END VDD
END NAND2XL

MACRO NAND2X4
    CLASS CORE ;
    FOREIGN NAND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.030 4.480 2.660 ;
        RECT  4.100 1.030 4.440 3.350 ;
        RECT  1.880 1.290 4.100 1.590 ;
        RECT  0.820 3.010 4.100 3.350 ;
        RECT  1.540 1.190 1.880 1.590 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.000 2.420 3.055 2.760 ;
        RECT  2.715 2.420 3.000 2.780 ;
        RECT  1.105 2.550 2.715 2.780 ;
        RECT  0.655 2.405 1.105 2.780 ;
        RECT  0.600 2.405 0.655 2.745 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.640 1.960 3.870 2.740 ;
        RECT  3.440 1.960 3.640 2.405 ;
        RECT  2.470 1.960 3.440 2.190 ;
        RECT  2.150 1.845 2.470 2.190 ;
        RECT  1.870 1.960 2.150 2.190 ;
        RECT  1.585 1.960 1.870 2.320 ;
        RECT  1.530 1.980 1.585 2.320 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 -0.400 4.620 0.400 ;
        RECT  2.820 -0.400 3.160 1.060 ;
        RECT  0.620 -0.400 2.820 0.400 ;
        RECT  0.280 -0.400 0.620 0.575 ;
        RECT  0.000 -0.400 0.280 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.360 4.640 4.620 5.440 ;
        RECT  4.020 3.595 4.360 5.440 ;
        RECT  3.080 4.640 4.020 5.440 ;
        RECT  2.740 3.595 3.080 5.440 ;
        RECT  1.800 4.640 2.740 5.440 ;
        RECT  1.460 3.595 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.595 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NAND2X4

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.915 1.690 3.145 3.235 ;
        RECT  2.495 1.690 2.915 1.920 ;
        RECT  2.855 2.955 2.915 3.235 ;
        RECT  0.920 2.955 2.855 3.185 ;
        RECT  2.265 1.045 2.495 1.920 ;
        RECT  2.195 1.045 2.265 1.285 ;
        RECT  1.840 1.045 2.195 1.275 ;
        RECT  1.500 0.935 1.840 1.275 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.450 2.345 2.680 2.710 ;
        RECT  1.105 2.425 2.450 2.655 ;
        RECT  0.735 2.405 1.105 2.655 ;
        RECT  0.680 2.405 0.735 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.680 2.020 2.185 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 -0.400 3.300 0.400 ;
        RECT  2.780 -0.400 3.120 1.275 ;
        RECT  0.520 -0.400 2.780 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 4.640 3.300 5.440 ;
        RECT  0.770 4.465 3.120 5.440 ;
        RECT  0.000 4.640 0.770 5.440 ;
        END
    END VDD
END NAND2X2

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2XL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 1.260 1.860 3.120 ;
        RECT  1.630 1.185 1.800 3.120 ;
        RECT  1.460 1.185 1.630 1.540 ;
        RECT  1.160 2.890 1.630 3.120 ;
        RECT  0.820 2.890 1.160 3.230 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.840 0.520 2.510 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.225 1.390 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.400 1.980 0.400 ;
        RECT  0.180 -0.400 0.520 1.440 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 4.640 1.980 5.440 ;
        RECT  0.180 4.465 1.185 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END NAND2X1

MACRO MXI4XL
    CLASS CORE ;
    FOREIGN MXI4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.675 1.350 14.980 3.545 ;
        RECT  14.660 1.350 14.675 1.850 ;
        RECT  14.640 2.955 14.675 3.545 ;
        RECT  14.640 1.350 14.660 1.690 ;
        RECT  14.075 2.955 14.640 3.205 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 2.240 13.060 2.660 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 1.820 4.450 2.380 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 1.260 5.800 1.995 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.360 1.630 9.100 2.100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.595 1.285 3.745 1.515 ;
        RECT  3.365 1.285 3.595 2.050 ;
        RECT  3.230 1.710 3.365 2.050 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.020 0.730 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.100 -0.400 15.180 0.400 ;
        RECT  13.760 -0.400 14.100 0.575 ;
        RECT  12.380 -0.400 13.760 0.400 ;
        RECT  11.960 -0.400 12.380 0.915 ;
        RECT  8.860 -0.400 11.960 0.400 ;
        RECT  8.520 -0.400 8.860 0.575 ;
        RECT  5.550 -0.400 8.520 0.400 ;
        RECT  5.130 -0.400 5.550 0.985 ;
        RECT  3.830 -0.400 5.130 0.400 ;
        RECT  3.410 -0.400 3.830 0.985 ;
        RECT  0.800 -0.400 3.410 0.400 ;
        RECT  0.460 -0.400 0.800 0.575 ;
        RECT  0.000 -0.400 0.460 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 4.640 15.180 5.440 ;
        RECT  13.800 4.465 14.140 5.440 ;
        RECT  12.340 4.640 13.800 5.440 ;
        RECT  12.000 3.280 12.340 5.440 ;
        RECT  8.890 4.640 12.000 5.440 ;
        RECT  8.550 4.465 8.890 5.440 ;
        RECT  5.550 4.640 8.550 5.440 ;
        RECT  5.130 3.935 5.550 5.440 ;
        RECT  3.910 4.640 5.130 5.440 ;
        RECT  3.490 3.935 3.910 5.440 ;
        RECT  0.520 4.640 3.490 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.250 2.100 14.360 2.440 ;
        RECT  14.020 0.815 14.250 2.440 ;
        RECT  12.840 0.815 14.020 1.045 ;
        RECT  13.295 1.275 13.525 3.510 ;
        RECT  13.090 1.275 13.295 1.945 ;
        RECT  13.220 3.280 13.295 3.510 ;
        RECT  12.880 3.280 13.220 3.620 ;
        RECT  11.325 1.715 13.090 1.945 ;
        RECT  12.610 0.815 12.840 1.395 ;
        RECT  11.640 1.165 12.610 1.395 ;
        RECT  11.925 2.450 11.980 2.790 ;
        RECT  11.685 2.415 11.925 2.790 ;
        RECT  11.455 2.415 11.685 4.135 ;
        RECT  11.410 0.640 11.640 1.395 ;
        RECT  6.225 3.905 11.455 4.135 ;
        RECT  10.390 0.640 11.410 0.870 ;
        RECT  11.095 1.715 11.325 2.070 ;
        RECT  10.855 1.105 11.170 1.445 ;
        RECT  10.855 3.280 11.140 3.620 ;
        RECT  10.625 1.105 10.855 3.620 ;
        RECT  10.335 0.640 10.390 1.400 ;
        RECT  10.335 3.060 10.390 3.400 ;
        RECT  10.160 0.640 10.335 3.400 ;
        RECT  10.105 1.060 10.160 3.400 ;
        RECT  10.050 1.060 10.105 1.400 ;
        RECT  10.050 3.060 10.105 3.400 ;
        RECT  9.435 1.050 9.665 3.520 ;
        RECT  9.320 1.050 9.435 1.390 ;
        RECT  9.290 3.180 9.435 3.520 ;
        RECT  8.770 2.370 9.110 2.710 ;
        RECT  8.555 2.480 8.770 2.710 ;
        RECT  8.325 2.480 8.555 3.510 ;
        RECT  7.500 3.280 8.325 3.510 ;
        RECT  8.035 1.020 8.150 1.360 ;
        RECT  8.035 2.710 8.090 3.050 ;
        RECT  7.805 1.020 8.035 3.050 ;
        RECT  7.750 2.710 7.805 3.050 ;
        RECT  7.270 1.080 7.500 3.510 ;
        RECT  6.930 1.080 7.270 1.420 ;
        RECT  6.820 3.280 7.270 3.510 ;
        RECT  6.765 1.675 6.995 3.045 ;
        RECT  6.335 1.675 6.765 1.905 ;
        RECT  5.990 2.815 6.765 3.045 ;
        RECT  6.165 2.165 6.475 2.555 ;
        RECT  6.335 1.080 6.390 1.420 ;
        RECT  6.105 1.080 6.335 1.905 ;
        RECT  5.995 3.395 6.225 4.135 ;
        RECT  5.015 2.325 6.165 2.555 ;
        RECT  6.050 1.080 6.105 1.420 ;
        RECT  1.755 3.395 5.995 3.625 ;
        RECT  4.785 1.315 5.015 3.085 ;
        RECT  4.670 1.315 4.785 1.545 ;
        RECT  4.750 2.800 4.785 3.085 ;
        RECT  4.410 2.800 4.750 3.140 ;
        RECT  4.335 1.180 4.670 1.545 ;
        RECT  3.605 2.855 4.410 3.085 ;
        RECT  4.330 1.180 4.335 1.520 ;
        RECT  3.375 2.375 3.605 3.085 ;
        RECT  2.870 2.375 3.375 2.605 ;
        RECT  2.275 2.895 3.030 3.125 ;
        RECT  2.755 1.180 2.890 1.520 ;
        RECT  2.570 2.200 2.870 2.610 ;
        RECT  2.525 1.180 2.755 1.970 ;
        RECT  2.565 2.240 2.570 2.605 ;
        RECT  2.275 1.740 2.525 1.970 ;
        RECT  2.045 1.740 2.275 3.125 ;
        RECT  1.755 1.235 1.995 1.465 ;
        RECT  1.525 1.235 1.755 3.625 ;
        RECT  1.235 2.920 1.290 3.260 ;
        RECT  1.005 1.180 1.235 3.260 ;
        RECT  0.750 1.180 1.005 1.520 ;
        RECT  0.950 2.920 1.005 3.260 ;
    END
END MXI4XL

MACRO MXI4X4
    CLASS CORE ;
    FOREIGN MXI4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI4XL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.380 0.985 15.700 3.795 ;
        RECT  15.320 0.770 15.380 4.265 ;
        RECT  15.040 0.770 15.320 1.580 ;
        RECT  15.040 2.985 15.320 4.265 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.020 2.310 12.580 2.690 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.520 2.380 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.625 1.820 5.800 2.100 ;
        RECT  5.245 1.820 5.625 2.295 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.590 1.260 9.045 1.540 ;
        RECT  8.365 1.260 8.590 2.355 ;
        RECT  8.360 1.285 8.365 2.355 ;
        RECT  8.260 1.990 8.360 2.355 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 1.970 3.845 2.295 ;
        RECT  3.440 1.270 3.820 2.295 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.210 0.780 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.140 -0.400 16.500 0.400 ;
        RECT  15.800 -0.400 16.140 0.575 ;
        RECT  14.620 -0.400 15.800 0.400 ;
        RECT  14.280 -0.400 14.620 0.575 ;
        RECT  13.160 -0.400 14.280 0.400 ;
        RECT  12.820 -0.400 13.160 0.575 ;
        RECT  8.845 -0.400 12.820 0.400 ;
        RECT  8.505 -0.400 8.845 0.975 ;
        RECT  5.495 -0.400 8.505 0.400 ;
        RECT  5.155 -0.400 5.495 1.030 ;
        RECT  3.970 -0.400 5.155 0.400 ;
        RECT  3.630 -0.400 3.970 0.985 ;
        RECT  0.570 -0.400 3.630 0.400 ;
        RECT  0.230 -0.400 0.570 1.275 ;
        RECT  0.000 -0.400 0.230 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.140 4.640 16.500 5.440 ;
        RECT  15.800 4.465 16.140 5.440 ;
        RECT  14.620 4.640 15.800 5.440 ;
        RECT  14.280 4.465 14.620 5.440 ;
        RECT  12.980 4.640 14.280 5.440 ;
        RECT  12.640 4.465 12.980 5.440 ;
        RECT  8.845 4.640 12.640 5.440 ;
        RECT  8.505 4.465 8.845 5.440 ;
        RECT  5.485 4.640 8.505 5.440 ;
        RECT  5.145 4.130 5.485 5.440 ;
        RECT  3.970 4.640 5.145 5.440 ;
        RECT  3.630 4.130 3.970 5.440 ;
        RECT  0.570 4.640 3.630 5.440 ;
        RECT  0.230 3.575 0.570 5.440 ;
        RECT  0.000 4.640 0.230 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.790 2.085 14.900 2.425 ;
        RECT  14.560 0.830 14.790 2.425 ;
        RECT  12.430 0.830 14.560 1.060 ;
        RECT  14.005 2.270 14.235 4.235 ;
        RECT  13.860 2.270 14.005 2.500 ;
        RECT  6.205 4.005 14.005 4.235 ;
        RECT  13.215 1.315 13.920 1.545 ;
        RECT  13.520 2.160 13.860 2.500 ;
        RECT  13.215 2.960 13.760 3.770 ;
        RECT  12.985 1.315 13.215 3.770 ;
        RECT  11.205 3.540 12.985 3.770 ;
        RECT  12.200 0.685 12.430 1.060 ;
        RECT  11.790 1.420 12.215 1.650 ;
        RECT  10.385 0.685 12.200 0.915 ;
        RECT  11.790 3.080 12.180 3.310 ;
        RECT  11.560 1.420 11.790 3.310 ;
        RECT  11.010 3.345 11.205 3.770 ;
        RECT  11.010 1.535 11.060 1.900 ;
        RECT  10.780 1.535 11.010 3.770 ;
        RECT  10.330 3.345 10.430 3.685 ;
        RECT  10.330 0.685 10.385 1.330 ;
        RECT  10.155 0.685 10.330 3.685 ;
        RECT  10.100 0.990 10.155 3.685 ;
        RECT  10.045 0.990 10.100 1.330 ;
        RECT  9.480 0.745 9.710 3.680 ;
        RECT  9.245 0.745 9.480 0.975 ;
        RECT  9.000 2.080 9.230 3.770 ;
        RECT  7.285 3.540 9.000 3.770 ;
        RECT  7.530 1.425 7.760 3.085 ;
        RECT  7.055 0.740 7.285 3.770 ;
        RECT  6.630 0.740 7.055 0.970 ;
        RECT  6.595 3.540 7.055 3.770 ;
        RECT  6.585 1.360 6.815 3.215 ;
        RECT  5.925 1.360 6.585 1.590 ;
        RECT  5.835 2.985 6.585 3.215 ;
        RECT  5.980 2.320 6.355 2.755 ;
        RECT  5.975 3.670 6.205 4.235 ;
        RECT  4.980 2.525 5.980 2.755 ;
        RECT  2.245 3.670 5.975 3.900 ;
        RECT  4.750 1.245 4.980 3.125 ;
        RECT  4.410 1.245 4.750 1.585 ;
        RECT  3.820 2.895 4.750 3.125 ;
        RECT  3.590 2.525 3.820 3.125 ;
        RECT  3.090 2.525 3.590 2.755 ;
        RECT  2.630 2.985 3.230 3.215 ;
        RECT  2.940 1.440 3.210 1.820 ;
        RECT  2.860 2.210 3.090 2.755 ;
        RECT  2.630 1.590 2.940 1.820 ;
        RECT  2.400 1.590 2.630 3.215 ;
        RECT  2.135 0.935 2.450 1.275 ;
        RECT  2.135 3.560 2.245 3.900 ;
        RECT  1.905 0.935 2.135 3.900 ;
        RECT  1.240 0.950 1.450 1.790 ;
        RECT  1.010 0.950 1.240 3.090 ;
    END
END MXI4X4

MACRO MXI4X2
    CLASS CORE ;
    FOREIGN MXI4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI4XL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.415 0.770 15.645 4.230 ;
        RECT  15.280 0.770 15.415 1.580 ;
        RECT  15.395 2.635 15.415 4.230 ;
        RECT  15.270 2.795 15.395 4.230 ;
        RECT  14.660 2.795 15.270 3.220 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.020 1.820 12.715 2.200 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 1.820 4.480 2.380 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 1.270 5.840 2.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.645 1.260 9.100 1.540 ;
        RECT  8.420 1.260 8.645 2.355 ;
        RECT  8.415 1.285 8.420 2.355 ;
        RECT  8.315 1.990 8.415 2.355 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.655 1.285 3.745 1.515 ;
        RECT  3.425 1.285 3.655 2.215 ;
        RECT  3.250 1.890 3.425 2.215 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.210 0.790 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.800 -0.400 15.840 0.400 ;
        RECT  14.460 -0.400 14.800 0.575 ;
        RECT  13.080 -0.400 14.460 0.400 ;
        RECT  12.740 -0.400 13.080 0.575 ;
        RECT  8.900 -0.400 12.740 0.400 ;
        RECT  8.560 -0.400 8.900 0.975 ;
        RECT  5.740 -0.400 8.560 0.400 ;
        RECT  5.400 -0.400 5.740 0.975 ;
        RECT  3.930 -0.400 5.400 0.400 ;
        RECT  3.590 -0.400 3.930 0.985 ;
        RECT  0.570 -0.400 3.590 0.400 ;
        RECT  0.230 -0.400 0.570 1.445 ;
        RECT  0.000 -0.400 0.230 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.710 4.640 15.840 5.440 ;
        RECT  14.370 4.465 14.710 5.440 ;
        RECT  12.950 4.640 14.370 5.440 ;
        RECT  12.610 4.465 12.950 5.440 ;
        RECT  8.900 4.640 12.610 5.440 ;
        RECT  8.560 4.465 8.900 5.440 ;
        RECT  5.540 4.640 8.560 5.440 ;
        RECT  5.200 3.945 5.540 5.440 ;
        RECT  3.930 4.640 5.200 5.440 ;
        RECT  3.590 3.945 3.930 5.440 ;
        RECT  0.570 4.640 3.590 5.440 ;
        RECT  0.230 3.065 0.570 5.440 ;
        RECT  0.000 4.640 0.230 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.990 2.085 15.100 2.425 ;
        RECT  14.760 0.830 14.990 2.425 ;
        RECT  12.485 0.830 14.760 1.060 ;
        RECT  14.015 2.275 14.245 4.235 ;
        RECT  13.235 1.315 14.020 1.545 ;
        RECT  13.880 2.275 14.015 2.505 ;
        RECT  6.205 4.005 14.015 4.235 ;
        RECT  13.595 2.160 13.880 2.505 ;
        RECT  13.235 3.195 13.725 3.585 ;
        RECT  13.540 2.160 13.595 2.500 ;
        RECT  13.005 1.315 13.235 3.585 ;
        RECT  11.260 3.355 13.005 3.585 ;
        RECT  12.255 0.685 12.485 1.060 ;
        RECT  11.980 2.675 12.345 3.085 ;
        RECT  10.440 0.685 12.255 0.915 ;
        RECT  11.715 2.675 11.980 2.905 ;
        RECT  11.715 1.315 11.940 1.545 ;
        RECT  11.485 1.315 11.715 2.905 ;
        RECT  11.355 1.870 11.485 2.290 ;
        RECT  11.065 3.220 11.260 3.585 ;
        RECT  11.065 1.205 11.145 1.570 ;
        RECT  10.835 1.205 11.065 3.585 ;
        RECT  10.385 3.345 10.485 3.685 ;
        RECT  10.385 0.685 10.440 1.440 ;
        RECT  10.210 0.685 10.385 3.685 ;
        RECT  10.155 1.100 10.210 3.685 ;
        RECT  10.100 1.100 10.155 1.440 ;
        RECT  9.535 0.745 9.765 3.685 ;
        RECT  9.340 0.745 9.535 0.975 ;
        RECT  9.055 2.080 9.285 3.770 ;
        RECT  7.505 3.540 9.055 3.770 ;
        RECT  7.795 1.060 8.025 3.260 ;
        RECT  7.275 1.060 7.505 3.770 ;
        RECT  6.980 1.060 7.275 1.400 ;
        RECT  6.740 3.540 7.275 3.770 ;
        RECT  6.755 1.830 6.985 3.250 ;
        RECT  6.560 1.830 6.755 2.060 ;
        RECT  5.980 3.020 6.755 3.250 ;
        RECT  6.330 1.060 6.560 2.060 ;
        RECT  6.235 2.295 6.465 2.790 ;
        RECT  6.220 1.060 6.330 1.400 ;
        RECT  5.015 2.560 6.235 2.790 ;
        RECT  5.975 3.485 6.205 4.235 ;
        RECT  1.815 3.485 5.975 3.715 ;
        RECT  4.785 1.205 5.015 3.125 ;
        RECT  4.410 1.205 4.785 1.435 ;
        RECT  3.495 2.895 4.785 3.125 ;
        RECT  3.265 2.500 3.495 3.125 ;
        RECT  2.855 2.500 3.265 2.730 ;
        RECT  2.910 1.090 3.020 1.430 ;
        RECT  2.335 2.960 2.950 3.190 ;
        RECT  2.680 1.090 2.910 1.845 ;
        RECT  2.625 2.140 2.855 2.730 ;
        RECT  2.335 1.615 2.680 1.845 ;
        RECT  2.105 1.615 2.335 3.190 ;
        RECT  1.815 0.995 2.150 1.335 ;
        RECT  1.585 0.995 1.815 3.715 ;
        RECT  1.065 1.105 1.295 3.430 ;
    END
END MXI4X2

MACRO MXI4X1
    CLASS CORE ;
    FOREIGN MXI4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI4XL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.675 1.350 14.980 3.785 ;
        RECT  14.660 1.350 14.675 1.850 ;
        RECT  14.640 2.955 14.675 3.785 ;
        RECT  14.640 1.350 14.660 1.690 ;
        RECT  14.075 2.955 14.640 3.205 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 2.240 13.060 2.660 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 1.820 4.450 2.380 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 1.260 5.830 1.830 ;
        RECT  5.735 1.260 5.790 1.970 ;
        RECT  5.495 1.260 5.735 1.995 ;
        RECT  5.450 1.260 5.495 1.970 ;
        RECT  5.410 1.260 5.450 1.830 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.360 1.630 9.100 2.100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.595 1.285 3.745 1.515 ;
        RECT  3.365 1.285 3.595 2.050 ;
        RECT  3.230 1.710 3.365 2.050 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.020 0.730 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.100 -0.400 15.180 0.400 ;
        RECT  13.760 -0.400 14.100 0.575 ;
        RECT  12.380 -0.400 13.760 0.400 ;
        RECT  11.960 -0.400 12.380 0.915 ;
        RECT  8.860 -0.400 11.960 0.400 ;
        RECT  8.520 -0.400 8.860 0.575 ;
        RECT  5.550 -0.400 8.520 0.400 ;
        RECT  5.130 -0.400 5.550 0.985 ;
        RECT  3.830 -0.400 5.130 0.400 ;
        RECT  3.410 -0.400 3.830 0.985 ;
        RECT  0.800 -0.400 3.410 0.400 ;
        RECT  0.460 -0.400 0.800 0.575 ;
        RECT  0.000 -0.400 0.460 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 4.640 15.180 5.440 ;
        RECT  13.800 4.465 14.140 5.440 ;
        RECT  12.340 4.640 13.800 5.440 ;
        RECT  12.000 3.290 12.340 5.440 ;
        RECT  8.890 4.640 12.000 5.440 ;
        RECT  8.550 4.465 8.890 5.440 ;
        RECT  5.550 4.640 8.550 5.440 ;
        RECT  5.130 3.935 5.550 5.440 ;
        RECT  3.910 4.640 5.130 5.440 ;
        RECT  3.490 3.935 3.910 5.440 ;
        RECT  0.520 4.640 3.490 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.250 2.100 14.360 2.440 ;
        RECT  14.020 0.815 14.250 2.440 ;
        RECT  12.845 0.815 14.020 1.045 ;
        RECT  13.295 1.290 13.525 3.240 ;
        RECT  13.090 1.290 13.295 1.945 ;
        RECT  13.220 3.010 13.295 3.240 ;
        RECT  12.880 3.010 13.220 3.350 ;
        RECT  11.325 1.715 13.090 1.945 ;
        RECT  12.615 0.815 12.845 1.395 ;
        RECT  11.640 1.165 12.615 1.395 ;
        RECT  11.925 2.450 11.980 2.790 ;
        RECT  11.685 2.415 11.925 2.790 ;
        RECT  11.455 2.415 11.685 4.135 ;
        RECT  11.410 0.640 11.640 1.395 ;
        RECT  6.225 3.905 11.455 4.135 ;
        RECT  10.335 0.640 11.410 0.870 ;
        RECT  11.095 1.715 11.325 2.070 ;
        RECT  10.855 1.160 11.170 1.390 ;
        RECT  10.855 3.060 11.140 3.400 ;
        RECT  10.625 1.160 10.855 3.400 ;
        RECT  10.105 0.640 10.335 3.425 ;
        RECT  9.435 1.025 9.665 3.400 ;
        RECT  9.345 1.025 9.435 1.390 ;
        RECT  9.270 3.060 9.435 3.400 ;
        RECT  9.290 1.050 9.345 1.390 ;
        RECT  8.555 2.425 9.110 2.655 ;
        RECT  8.325 2.425 8.555 3.595 ;
        RECT  7.515 3.365 8.325 3.595 ;
        RECT  8.035 1.030 8.095 1.420 ;
        RECT  7.805 1.030 8.035 3.050 ;
        RECT  7.285 1.110 7.515 3.595 ;
        RECT  7.270 1.110 7.285 1.340 ;
        RECT  6.820 3.365 7.285 3.595 ;
        RECT  6.930 1.000 7.270 1.340 ;
        RECT  6.765 1.645 6.995 3.075 ;
        RECT  6.335 1.645 6.765 1.875 ;
        RECT  5.990 2.845 6.765 3.075 ;
        RECT  6.165 2.165 6.475 2.555 ;
        RECT  6.105 1.080 6.335 1.875 ;
        RECT  5.995 3.415 6.225 4.135 ;
        RECT  5.015 2.325 6.165 2.555 ;
        RECT  1.755 3.415 5.995 3.645 ;
        RECT  4.785 1.315 5.015 3.085 ;
        RECT  4.670 1.315 4.785 1.545 ;
        RECT  3.605 2.855 4.785 3.085 ;
        RECT  4.335 1.180 4.670 1.545 ;
        RECT  4.330 1.180 4.335 1.520 ;
        RECT  3.375 2.375 3.605 3.085 ;
        RECT  2.870 2.375 3.375 2.605 ;
        RECT  2.275 2.895 3.030 3.125 ;
        RECT  2.755 1.180 2.890 1.520 ;
        RECT  2.570 2.200 2.870 2.610 ;
        RECT  2.525 1.180 2.755 1.925 ;
        RECT  2.565 2.240 2.570 2.605 ;
        RECT  2.275 1.695 2.525 1.925 ;
        RECT  2.045 1.695 2.275 3.125 ;
        RECT  1.755 1.235 1.995 1.465 ;
        RECT  1.525 1.235 1.755 3.645 ;
        RECT  1.005 1.155 1.235 3.300 ;
        RECT  0.805 1.155 1.005 1.520 ;
        RECT  0.750 1.180 0.805 1.520 ;
    END
END MXI4X1

MACRO MXI2XL
    CLASS CORE ;
    FOREIGN MXI2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 2.405 3.085 3.440 ;
        RECT  2.945 1.180 3.000 1.520 ;
        RECT  2.715 1.180 2.945 3.440 ;
        RECT  2.660 1.180 2.715 1.520 ;
        RECT  2.660 3.100 2.715 3.440 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.705 2.200 1.180 2.660 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.820 1.880 2.330 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.820 4.480 2.280 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.430 -0.400 4.620 0.400 ;
        RECT  4.090 -0.400 4.430 0.575 ;
        RECT  1.435 -0.400 4.090 0.400 ;
        RECT  1.095 -0.400 1.435 1.520 ;
        RECT  0.000 -0.400 1.095 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.445 4.640 4.620 5.440 ;
        RECT  4.095 4.405 4.445 5.440 ;
        RECT  1.420 4.640 4.095 5.440 ;
        RECT  1.080 3.890 1.420 5.440 ;
        RECT  0.000 4.640 1.080 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.695 3.100 3.800 3.440 ;
        RECT  3.695 1.170 3.760 1.510 ;
        RECT  3.465 1.170 3.695 3.440 ;
        RECT  3.420 1.170 3.465 1.510 ;
        RECT  3.460 3.100 3.465 3.440 ;
        RECT  2.325 3.905 2.480 4.245 ;
        RECT  2.175 1.180 2.405 3.190 ;
        RECT  2.095 3.425 2.325 4.245 ;
        RECT  1.900 1.180 2.175 1.520 ;
        RECT  1.880 2.850 2.175 3.190 ;
        RECT  0.540 3.425 2.095 3.655 ;
        RECT  0.405 1.180 0.580 1.520 ;
        RECT  0.405 3.270 0.540 3.655 ;
        RECT  0.175 1.180 0.405 3.655 ;
    END
END MXI2XL

MACRO MXI2X4
    CLASS CORE ;
    FOREIGN MXI2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI2XL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.610 0.720 5.930 1.100 ;
        RECT  4.270 3.585 5.645 3.815 ;
        RECT  4.490 0.720 5.610 0.950 ;
        RECT  4.480 0.720 4.490 1.070 ;
        RECT  4.270 0.700 4.480 2.100 ;
        RECT  4.100 0.700 4.270 3.815 ;
        RECT  3.060 0.720 4.100 0.950 ;
        RECT  4.040 1.845 4.100 3.815 ;
        RECT  3.745 3.500 4.040 3.815 ;
        RECT  2.565 3.585 3.745 3.815 ;
        RECT  2.720 0.720 3.060 1.060 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.920 4.005 6.260 4.345 ;
        RECT  5.420 4.060 5.920 4.345 ;
        RECT  2.315 4.115 5.420 4.345 ;
        RECT  2.085 3.960 2.315 4.345 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.400 2.160 8.090 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.210 1.500 2.550 ;
        RECT  0.875 2.210 1.105 2.635 ;
        RECT  0.560 2.210 0.875 2.550 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.060 -0.400 9.240 0.400 ;
        RECT  8.720 -0.400 9.060 1.050 ;
        RECT  7.680 -0.400 8.720 0.400 ;
        RECT  7.340 -0.400 7.680 0.575 ;
        RECT  1.845 -0.400 7.340 0.400 ;
        RECT  1.505 -0.400 1.845 1.050 ;
        RECT  0.540 -0.400 1.505 0.400 ;
        RECT  0.200 -0.400 0.540 1.070 ;
        RECT  0.000 -0.400 0.200 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.060 4.640 9.240 5.440 ;
        RECT  8.720 4.050 9.060 5.440 ;
        RECT  7.655 4.640 8.720 5.440 ;
        RECT  7.315 3.700 7.655 5.440 ;
        RECT  1.785 4.640 7.315 5.440 ;
        RECT  1.555 4.050 1.785 5.440 ;
        RECT  0.540 4.640 1.555 5.440 ;
        RECT  0.200 4.060 0.540 5.440 ;
        RECT  0.000 4.640 0.200 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.665 1.525 8.895 3.190 ;
        RECT  8.400 1.525 8.665 1.755 ;
        RECT  8.395 2.960 8.665 3.190 ;
        RECT  8.285 1.410 8.400 1.755 ;
        RECT  8.055 2.960 8.395 3.635 ;
        RECT  8.115 0.930 8.285 1.755 ;
        RECT  8.060 0.930 8.115 1.750 ;
        RECT  8.055 0.930 8.060 1.695 ;
        RECT  6.395 0.930 8.055 1.160 ;
        RECT  6.855 2.780 6.995 3.210 ;
        RECT  6.625 1.410 6.855 3.210 ;
        RECT  6.260 2.980 6.625 3.210 ;
        RECT  6.165 0.930 6.395 1.695 ;
        RECT  5.920 2.980 6.260 3.320 ;
        RECT  5.180 1.465 6.165 1.695 ;
        RECT  4.950 1.465 5.180 3.080 ;
        RECT  4.935 2.850 4.950 3.080 ;
        RECT  4.595 2.850 4.935 3.190 ;
        RECT  3.355 1.410 3.695 1.750 ;
        RECT  3.230 2.760 3.570 3.155 ;
        RECT  3.235 1.520 3.355 1.750 ;
        RECT  3.005 1.520 3.235 1.885 ;
        RECT  2.075 2.925 3.230 3.155 ;
        RECT  2.075 1.655 3.005 1.885 ;
        RECT  1.845 1.655 2.075 3.165 ;
        RECT  1.200 1.655 1.845 1.885 ;
        RECT  1.200 2.925 1.845 3.165 ;
        RECT  0.860 1.410 1.200 1.885 ;
        RECT  0.915 2.925 1.200 3.300 ;
        RECT  0.860 2.935 0.915 3.300 ;
    END
END MXI2X4

MACRO MXI2X2
    CLASS CORE ;
    FOREIGN MXI2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.330 1.230 3.560 3.730 ;
        RECT  3.160 3.500 3.330 3.730 ;
        RECT  2.700 3.500 3.160 4.220 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.675 2.755 1.180 3.220 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.125 1.860 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.720 1.820 5.140 2.420 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 -0.400 5.280 0.400 ;
        RECT  4.760 -0.400 5.100 0.575 ;
        RECT  1.730 -0.400 4.760 0.400 ;
        RECT  1.390 -0.400 1.730 1.160 ;
        RECT  0.000 -0.400 1.390 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 4.640 5.280 5.440 ;
        RECT  4.760 3.115 5.100 5.440 ;
        RECT  1.420 4.640 4.760 5.440 ;
        RECT  1.080 3.520 1.420 5.440 ;
        RECT  0.000 4.640 1.080 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.255 1.410 4.485 3.320 ;
        RECT  4.205 3.090 4.255 3.320 ;
        RECT  3.865 3.090 4.205 4.030 ;
        RECT  3.790 0.685 4.020 2.400 ;
        RECT  2.320 0.685 3.790 0.915 ;
        RECT  2.870 1.370 3.100 3.205 ;
        RECT  2.555 1.370 2.870 1.710 ;
        RECT  2.200 2.975 2.870 3.205 ;
        RECT  2.320 2.170 2.625 2.550 ;
        RECT  2.090 0.685 2.320 2.550 ;
        RECT  1.860 2.975 2.200 4.255 ;
        RECT  0.970 1.625 2.090 1.855 ;
        RECT  0.740 1.080 0.970 1.855 ;
        RECT  0.630 1.080 0.740 1.460 ;
        RECT  0.410 1.230 0.630 1.460 ;
        RECT  0.410 3.510 0.520 3.850 ;
        RECT  0.180 1.230 0.410 3.850 ;
    END
END MXI2X2

MACRO MXI2X1
    CLASS CORE ;
    FOREIGN MXI2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 2.405 3.085 3.380 ;
        RECT  2.945 1.180 3.000 1.520 ;
        RECT  2.715 1.180 2.945 3.380 ;
        RECT  2.660 1.180 2.715 1.520 ;
        RECT  2.660 3.040 2.715 3.380 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.705 2.200 1.180 2.660 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.820 1.880 2.330 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.820 4.480 2.280 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.430 -0.400 4.620 0.400 ;
        RECT  4.090 -0.400 4.430 0.575 ;
        RECT  1.460 -0.400 4.090 0.400 ;
        RECT  1.120 -0.400 1.460 1.520 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.445 4.640 4.620 5.440 ;
        RECT  4.095 4.405 4.445 5.440 ;
        RECT  1.420 4.640 4.095 5.440 ;
        RECT  1.080 3.945 1.420 5.440 ;
        RECT  0.000 4.640 1.080 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.695 2.980 3.800 3.320 ;
        RECT  3.695 1.170 3.760 1.510 ;
        RECT  3.465 1.170 3.695 3.320 ;
        RECT  3.420 1.170 3.465 1.510 ;
        RECT  3.460 2.980 3.465 3.320 ;
        RECT  2.325 3.920 2.480 4.260 ;
        RECT  2.175 1.180 2.405 3.190 ;
        RECT  2.095 3.425 2.325 4.260 ;
        RECT  1.900 1.180 2.175 1.520 ;
        RECT  1.880 2.850 2.175 3.190 ;
        RECT  0.540 3.425 2.095 3.655 ;
        RECT  0.580 1.225 0.585 1.545 ;
        RECT  0.405 1.225 0.580 1.600 ;
        RECT  0.405 3.090 0.540 3.655 ;
        RECT  0.175 1.225 0.405 3.655 ;
    END
END MXI2X1

MACRO MX4XL
    CLASS CORE ;
    FOREIGN MX4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.705 1.280 12.990 4.170 ;
        RECT  12.650 1.280 12.705 1.850 ;
        RECT  12.650 3.750 12.705 4.170 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 0.640 9.760 0.980 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.050 2.360 4.545 2.780 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 1.820 3.820 2.255 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 1.930 0.770 2.270 ;
        RECT  0.140 1.820 0.520 2.270 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.280 1.815 5.890 2.185 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 1.820 8.565 2.450 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.230 -0.400 13.200 0.400 ;
        RECT  11.890 -0.400 12.230 0.575 ;
        RECT  8.730 -0.400 11.890 0.400 ;
        RECT  8.390 -0.400 8.730 0.575 ;
        RECT  5.460 -0.400 8.390 0.400 ;
        RECT  5.120 -0.400 5.460 1.440 ;
        RECT  3.795 -0.400 5.120 0.400 ;
        RECT  3.455 -0.400 3.795 1.440 ;
        RECT  0.540 -0.400 3.455 0.400 ;
        RECT  0.200 -0.400 0.540 0.575 ;
        RECT  0.000 -0.400 0.200 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.210 4.640 13.200 5.440 ;
        RECT  11.870 4.465 12.210 5.440 ;
        RECT  8.730 4.640 11.870 5.440 ;
        RECT  8.390 4.465 8.730 5.440 ;
        RECT  5.480 4.640 8.390 5.440 ;
        RECT  5.140 3.960 5.480 5.440 ;
        RECT  3.790 4.640 5.140 5.440 ;
        RECT  3.450 3.960 3.790 5.440 ;
        RECT  0.540 4.640 3.450 5.440 ;
        RECT  0.200 4.465 0.540 5.440 ;
        RECT  0.000 4.640 0.200 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.165 2.020 12.435 2.370 ;
        RECT  11.935 0.860 12.165 2.370 ;
        RECT  11.915 2.880 11.960 3.220 ;
        RECT  10.950 0.860 11.935 1.090 ;
        RECT  11.685 2.880 11.915 4.235 ;
        RECT  11.615 2.880 11.685 3.220 ;
        RECT  6.340 4.005 11.685 4.235 ;
        RECT  11.385 1.370 11.615 3.220 ;
        RECT  10.950 3.285 11.150 3.625 ;
        RECT  10.720 0.860 10.950 3.625 ;
        RECT  10.565 1.305 10.720 1.645 ;
        RECT  10.280 3.370 10.390 3.765 ;
        RECT  10.050 1.305 10.280 3.765 ;
        RECT  9.815 1.305 10.050 1.645 ;
        RECT  7.340 3.535 10.050 3.765 ;
        RECT  9.440 1.920 9.550 3.250 ;
        RECT  9.320 1.300 9.440 3.250 ;
        RECT  9.210 1.300 9.320 2.260 ;
        RECT  9.210 2.910 9.320 3.250 ;
        RECT  9.100 1.300 9.210 1.640 ;
        RECT  7.825 2.910 8.060 3.250 ;
        RECT  7.595 1.180 7.825 3.250 ;
        RECT  7.120 1.210 7.340 3.765 ;
        RECT  7.110 1.130 7.120 3.765 ;
        RECT  6.780 1.130 7.110 1.470 ;
        RECT  6.900 3.535 7.110 3.765 ;
        RECT  6.650 1.725 6.880 3.265 ;
        RECT  6.490 1.725 6.650 1.955 ;
        RECT  6.055 3.035 6.650 3.265 ;
        RECT  6.330 1.210 6.490 1.955 ;
        RECT  6.140 2.300 6.420 2.675 ;
        RECT  6.110 3.495 6.340 4.235 ;
        RECT  6.260 1.100 6.330 1.955 ;
        RECT  5.990 1.100 6.260 1.440 ;
        RECT  5.035 2.425 6.140 2.675 ;
        RECT  2.170 3.495 6.110 3.725 ;
        RECT  4.805 1.870 5.035 3.265 ;
        RECT  4.670 1.870 4.805 2.100 ;
        RECT  3.565 3.035 4.805 3.265 ;
        RECT  4.330 1.240 4.670 2.100 ;
        RECT  3.335 2.505 3.565 3.265 ;
        RECT  2.755 2.505 3.335 2.735 ;
        RECT  2.245 3.035 2.990 3.265 ;
        RECT  2.840 1.100 2.950 1.440 ;
        RECT  2.610 1.100 2.840 2.005 ;
        RECT  2.475 2.280 2.755 2.735 ;
        RECT  2.245 1.775 2.610 2.005 ;
        RECT  2.015 1.775 2.245 3.265 ;
        RECT  1.830 1.100 2.170 1.440 ;
        RECT  1.830 3.495 2.170 3.835 ;
        RECT  1.780 1.170 1.830 1.440 ;
        RECT  1.780 3.495 1.830 3.725 ;
        RECT  1.550 1.170 1.780 3.725 ;
        RECT  1.090 1.100 1.320 3.415 ;
    END
END MX4XL

MACRO MX4X4
    CLASS CORE ;
    FOREIGN MX4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX4XL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.660 1.345 15.040 3.780 ;
        RECT  14.575 1.345 14.660 1.780 ;
        RECT  14.575 2.760 14.660 3.780 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.935 2.430 13.250 2.770 ;
        RECT  12.705 2.430 12.935 3.755 ;
        RECT  11.080 3.525 12.705 3.755 ;
        RECT  10.700 3.525 11.080 3.860 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.635 3.995 7.865 4.340 ;
        RECT  2.855 3.995 7.635 4.225 ;
        RECT  2.425 3.995 2.855 4.260 ;
        RECT  2.375 3.995 2.425 4.315 ;
        RECT  2.330 4.030 2.375 4.315 ;
        RECT  1.990 4.030 2.330 4.370 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 2.355 4.405 2.635 ;
        RECT  3.810 2.355 4.175 2.585 ;
        RECT  3.580 2.200 3.810 2.585 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.820 0.760 2.310 ;
        RECT  0.140 1.820 0.420 2.305 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.960 1.820 6.460 2.270 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.250 2.205 9.760 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.570 -0.400 15.840 0.400 ;
        RECT  15.230 -0.400 15.570 1.080 ;
        RECT  14.250 -0.400 15.230 0.400 ;
        RECT  13.910 -0.400 14.250 1.005 ;
        RECT  9.835 -0.400 13.910 0.400 ;
        RECT  9.495 -0.400 9.835 0.575 ;
        RECT  6.070 -0.400 9.495 0.400 ;
        RECT  5.730 -0.400 6.070 0.575 ;
        RECT  4.320 -0.400 5.730 0.400 ;
        RECT  3.980 -0.400 4.320 0.575 ;
        RECT  0.520 -0.400 3.980 0.400 ;
        RECT  0.180 -0.400 0.520 1.590 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.570 4.640 15.840 5.440 ;
        RECT  15.230 4.060 15.570 5.440 ;
        RECT  14.250 4.640 15.230 5.440 ;
        RECT  13.910 4.060 14.250 5.440 ;
        RECT  9.830 4.640 13.910 5.440 ;
        RECT  9.490 4.465 9.830 5.440 ;
        RECT  6.070 4.640 9.490 5.440 ;
        RECT  5.730 4.465 6.070 5.440 ;
        RECT  4.195 4.640 5.730 5.440 ;
        RECT  3.855 4.465 4.195 5.440 ;
        RECT  0.520 4.640 3.855 5.440 ;
        RECT  0.180 3.115 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.885 1.255 14.115 3.305 ;
        RECT  13.345 1.255 13.885 1.485 ;
        RECT  13.405 3.075 13.885 3.305 ;
        RECT  13.310 1.715 13.635 2.135 ;
        RECT  13.175 3.075 13.405 4.375 ;
        RECT  13.005 0.660 13.345 1.485 ;
        RECT  12.510 1.835 13.310 2.065 ;
        RECT  10.350 4.145 13.175 4.375 ;
        RECT  12.215 0.815 12.510 2.065 ;
        RECT  12.170 0.815 12.215 3.200 ;
        RECT  11.985 1.835 12.170 3.200 ;
        RECT  11.820 2.860 11.985 3.200 ;
        RECT  11.605 0.840 11.715 1.690 ;
        RECT  11.385 0.840 11.605 2.485 ;
        RECT  11.385 2.860 11.440 3.200 ;
        RECT  11.375 0.840 11.385 3.200 ;
        RECT  8.310 0.840 11.375 1.070 ;
        RECT  11.155 2.255 11.375 3.200 ;
        RECT  11.100 2.860 11.155 3.200 ;
        RECT  10.540 1.410 11.125 1.750 ;
        RECT  10.540 2.890 10.595 3.230 ;
        RECT  10.310 1.410 10.540 3.230 ;
        RECT  10.120 3.945 10.350 4.375 ;
        RECT  10.255 1.410 10.310 1.750 ;
        RECT  10.255 2.890 10.310 3.230 ;
        RECT  8.415 3.945 10.120 4.175 ;
        RECT  8.940 1.330 9.050 1.670 ;
        RECT  8.940 2.905 9.050 3.715 ;
        RECT  8.710 1.330 8.940 3.715 ;
        RECT  8.185 3.535 8.415 4.175 ;
        RECT  8.125 0.840 8.310 1.300 ;
        RECT  5.910 3.535 8.185 3.765 ;
        RECT  8.125 2.850 8.180 3.190 ;
        RECT  7.925 0.840 8.125 3.190 ;
        RECT  7.895 0.865 7.925 3.190 ;
        RECT  7.840 2.850 7.895 3.190 ;
        RECT  7.375 1.380 7.605 3.245 ;
        RECT  6.860 1.380 7.375 1.720 ;
        RECT  6.830 3.015 7.375 3.245 ;
        RECT  6.875 0.630 7.200 0.860 ;
        RECT  7.085 2.210 7.140 2.550 ;
        RECT  6.800 2.210 7.085 2.730 ;
        RECT  6.645 0.630 6.875 1.095 ;
        RECT  6.490 2.960 6.830 3.300 ;
        RECT  5.085 2.500 6.800 2.730 ;
        RECT  3.190 0.865 6.645 1.095 ;
        RECT  5.680 3.465 5.910 3.765 ;
        RECT  4.430 3.465 5.680 3.695 ;
        RECT  5.010 1.455 5.085 2.730 ;
        RECT  4.780 1.455 5.010 3.235 ;
        RECT  4.720 1.455 4.780 1.725 ;
        RECT  4.670 2.895 4.780 3.235 ;
        RECT  3.285 1.455 4.720 1.685 ;
        RECT  4.200 3.420 4.430 3.695 ;
        RECT  1.960 3.420 4.200 3.650 ;
        RECT  3.080 2.850 3.420 3.190 ;
        RECT  3.055 1.455 3.285 2.540 ;
        RECT  2.850 0.720 3.190 1.095 ;
        RECT  2.530 2.905 3.080 3.135 ;
        RECT  2.770 2.200 3.055 2.540 ;
        RECT  2.530 1.365 2.820 1.705 ;
        RECT  2.300 1.365 2.530 3.135 ;
        RECT  1.925 0.780 1.965 1.590 ;
        RECT  1.925 3.420 1.960 3.760 ;
        RECT  1.695 0.780 1.925 3.760 ;
        RECT  1.625 0.780 1.695 1.590 ;
        RECT  1.620 3.420 1.695 3.760 ;
        RECT  1.010 0.780 1.240 4.055 ;
        RECT  0.900 0.780 1.010 1.590 ;
        RECT  0.900 3.115 1.010 4.055 ;
    END
END MX4X4

MACRO MX4X2
    CLASS CORE ;
    FOREIGN MX4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX4XL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.825 2.965 14.965 3.195 ;
        RECT  14.595 0.755 14.825 4.225 ;
        RECT  14.485 0.755 14.595 1.565 ;
        RECT  14.485 2.945 14.595 4.225 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.935 2.430 13.250 2.770 ;
        RECT  12.705 2.430 12.935 3.755 ;
        RECT  11.080 3.525 12.705 3.755 ;
        RECT  10.700 3.525 11.080 3.860 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.635 3.995 7.865 4.340 ;
        RECT  2.855 3.995 7.635 4.225 ;
        RECT  2.425 3.995 2.855 4.260 ;
        RECT  2.375 3.995 2.425 4.315 ;
        RECT  2.330 4.030 2.375 4.315 ;
        RECT  1.990 4.030 2.330 4.370 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 2.355 4.405 2.635 ;
        RECT  3.810 2.355 4.175 2.585 ;
        RECT  3.580 2.200 3.810 2.585 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.820 0.760 2.310 ;
        RECT  0.140 1.820 0.420 2.305 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.960 1.820 6.460 2.270 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.250 2.205 9.760 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.045 -0.400 15.180 0.400 ;
        RECT  13.705 -0.400 14.045 0.945 ;
        RECT  9.835 -0.400 13.705 0.400 ;
        RECT  9.495 -0.400 9.835 0.575 ;
        RECT  6.070 -0.400 9.495 0.400 ;
        RECT  5.730 -0.400 6.070 0.575 ;
        RECT  4.320 -0.400 5.730 0.400 ;
        RECT  3.980 -0.400 4.320 0.575 ;
        RECT  0.520 -0.400 3.980 0.400 ;
        RECT  0.180 -0.400 0.520 1.590 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.045 4.640 15.180 5.440 ;
        RECT  13.705 3.620 14.045 5.440 ;
        RECT  9.830 4.640 13.705 5.440 ;
        RECT  9.490 4.465 9.830 5.440 ;
        RECT  6.070 4.640 9.490 5.440 ;
        RECT  5.730 4.465 6.070 5.440 ;
        RECT  4.195 4.640 5.730 5.440 ;
        RECT  3.855 4.465 4.195 5.440 ;
        RECT  0.520 4.640 3.855 5.440 ;
        RECT  0.180 3.115 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.885 1.240 14.115 3.305 ;
        RECT  13.345 1.240 13.885 1.470 ;
        RECT  13.405 3.075 13.885 3.305 ;
        RECT  13.310 1.715 13.635 2.135 ;
        RECT  13.175 3.075 13.405 4.375 ;
        RECT  13.005 0.660 13.345 1.470 ;
        RECT  12.510 1.835 13.310 2.065 ;
        RECT  10.350 4.145 13.175 4.375 ;
        RECT  12.170 0.815 12.510 2.065 ;
        RECT  12.160 1.835 12.170 2.065 ;
        RECT  11.930 1.835 12.160 3.200 ;
        RECT  11.820 2.860 11.930 3.200 ;
        RECT  11.605 0.840 11.715 1.690 ;
        RECT  11.385 0.840 11.605 2.485 ;
        RECT  11.385 2.860 11.440 3.200 ;
        RECT  11.375 0.840 11.385 3.200 ;
        RECT  8.310 0.840 11.375 1.070 ;
        RECT  11.155 2.255 11.375 3.200 ;
        RECT  11.100 2.860 11.155 3.200 ;
        RECT  10.540 1.410 11.125 1.750 ;
        RECT  10.540 2.890 10.595 3.230 ;
        RECT  10.310 1.410 10.540 3.230 ;
        RECT  10.120 3.945 10.350 4.375 ;
        RECT  10.255 1.410 10.310 1.750 ;
        RECT  10.255 2.890 10.310 3.230 ;
        RECT  8.415 3.945 10.120 4.175 ;
        RECT  8.940 1.330 9.050 1.670 ;
        RECT  8.940 2.905 9.050 3.715 ;
        RECT  8.710 1.330 8.940 3.715 ;
        RECT  8.185 3.535 8.415 4.175 ;
        RECT  8.125 0.840 8.310 1.300 ;
        RECT  5.910 3.535 8.185 3.765 ;
        RECT  8.125 2.850 8.180 3.190 ;
        RECT  7.925 0.840 8.125 3.190 ;
        RECT  7.895 0.865 7.925 3.190 ;
        RECT  7.840 2.850 7.895 3.190 ;
        RECT  7.375 1.380 7.605 3.245 ;
        RECT  6.860 1.380 7.375 1.720 ;
        RECT  6.830 3.015 7.375 3.245 ;
        RECT  6.875 0.630 7.200 0.860 ;
        RECT  7.085 2.210 7.140 2.550 ;
        RECT  6.800 2.210 7.085 2.730 ;
        RECT  6.645 0.630 6.875 1.095 ;
        RECT  6.490 2.960 6.830 3.300 ;
        RECT  5.085 2.500 6.800 2.730 ;
        RECT  3.190 0.865 6.645 1.095 ;
        RECT  5.680 3.465 5.910 3.765 ;
        RECT  4.430 3.465 5.680 3.695 ;
        RECT  5.010 1.455 5.085 2.730 ;
        RECT  4.780 1.455 5.010 3.235 ;
        RECT  4.720 1.455 4.780 1.725 ;
        RECT  4.670 2.895 4.780 3.235 ;
        RECT  3.285 1.455 4.720 1.685 ;
        RECT  4.200 3.420 4.430 3.695 ;
        RECT  1.960 3.420 4.200 3.650 ;
        RECT  3.080 2.850 3.420 3.190 ;
        RECT  3.055 1.455 3.285 2.540 ;
        RECT  2.850 0.720 3.190 1.095 ;
        RECT  2.530 2.905 3.080 3.135 ;
        RECT  2.770 2.200 3.055 2.540 ;
        RECT  2.530 1.365 2.820 1.705 ;
        RECT  2.300 1.365 2.530 3.135 ;
        RECT  1.925 0.780 1.965 1.590 ;
        RECT  1.925 3.420 1.960 3.760 ;
        RECT  1.695 0.780 1.925 3.760 ;
        RECT  1.625 0.780 1.695 1.590 ;
        RECT  1.620 3.420 1.695 3.760 ;
        RECT  1.010 0.780 1.240 4.055 ;
        RECT  0.900 0.780 1.010 1.590 ;
        RECT  0.900 3.115 1.010 4.055 ;
    END
END MX4X2

MACRO MX4X1
    CLASS CORE ;
    FOREIGN MX4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX4XL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.705 1.280 12.990 4.405 ;
        RECT  12.650 1.280 12.705 1.850 ;
        RECT  12.650 3.595 12.705 4.405 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 0.640 9.760 0.980 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.050 2.360 4.545 2.780 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 1.820 3.820 2.255 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 1.930 0.770 2.270 ;
        RECT  0.140 1.820 0.520 2.270 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.280 1.815 5.890 2.185 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 1.820 8.565 2.450 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.230 -0.400 13.200 0.400 ;
        RECT  11.890 -0.400 12.230 0.575 ;
        RECT  8.730 -0.400 11.890 0.400 ;
        RECT  8.390 -0.400 8.730 0.575 ;
        RECT  5.460 -0.400 8.390 0.400 ;
        RECT  5.120 -0.400 5.460 1.470 ;
        RECT  3.770 -0.400 5.120 0.400 ;
        RECT  3.430 -0.400 3.770 1.380 ;
        RECT  0.540 -0.400 3.430 0.400 ;
        RECT  0.200 -0.400 0.540 0.575 ;
        RECT  0.000 -0.400 0.200 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.210 4.640 13.200 5.440 ;
        RECT  11.870 4.465 12.210 5.440 ;
        RECT  8.730 4.640 11.870 5.440 ;
        RECT  8.390 4.465 8.730 5.440 ;
        RECT  5.480 4.640 8.390 5.440 ;
        RECT  5.140 3.960 5.480 5.440 ;
        RECT  3.790 4.640 5.140 5.440 ;
        RECT  3.450 3.960 3.790 5.440 ;
        RECT  0.540 4.640 3.450 5.440 ;
        RECT  0.200 4.465 0.540 5.440 ;
        RECT  0.000 4.640 0.200 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.165 2.020 12.435 2.370 ;
        RECT  11.935 0.860 12.165 2.370 ;
        RECT  11.915 2.880 11.960 3.220 ;
        RECT  10.950 0.860 11.935 1.090 ;
        RECT  11.685 2.880 11.915 4.235 ;
        RECT  11.615 2.880 11.685 3.220 ;
        RECT  6.340 4.005 11.685 4.235 ;
        RECT  11.385 1.370 11.615 3.220 ;
        RECT  10.950 3.285 11.150 3.625 ;
        RECT  10.720 0.860 10.950 3.625 ;
        RECT  10.565 1.220 10.720 1.560 ;
        RECT  10.280 3.370 10.390 3.765 ;
        RECT  10.050 1.220 10.280 3.765 ;
        RECT  9.815 1.220 10.050 1.560 ;
        RECT  7.340 3.535 10.050 3.765 ;
        RECT  9.440 1.920 9.550 3.250 ;
        RECT  9.320 1.320 9.440 3.250 ;
        RECT  9.210 1.320 9.320 2.260 ;
        RECT  9.210 2.910 9.320 3.250 ;
        RECT  9.100 1.320 9.210 1.660 ;
        RECT  7.825 2.910 8.060 3.250 ;
        RECT  7.595 1.180 7.825 3.250 ;
        RECT  7.120 1.210 7.340 3.765 ;
        RECT  7.110 1.130 7.120 3.765 ;
        RECT  6.780 1.130 7.110 1.470 ;
        RECT  6.900 3.535 7.110 3.765 ;
        RECT  6.650 1.725 6.880 3.265 ;
        RECT  6.490 1.725 6.650 1.955 ;
        RECT  6.140 3.035 6.650 3.265 ;
        RECT  6.310 1.210 6.490 1.955 ;
        RECT  6.140 2.300 6.420 2.675 ;
        RECT  6.110 3.495 6.340 4.235 ;
        RECT  6.260 1.130 6.310 1.955 ;
        RECT  5.970 1.130 6.260 1.470 ;
        RECT  5.035 2.425 6.140 2.675 ;
        RECT  2.170 3.495 6.110 3.725 ;
        RECT  4.805 1.870 5.035 3.265 ;
        RECT  4.650 1.870 4.805 2.100 ;
        RECT  3.565 3.035 4.805 3.265 ;
        RECT  4.310 1.240 4.650 2.100 ;
        RECT  3.335 2.505 3.565 3.265 ;
        RECT  2.755 2.505 3.335 2.735 ;
        RECT  2.245 3.035 3.010 3.265 ;
        RECT  2.840 1.040 2.950 1.380 ;
        RECT  2.610 1.040 2.840 2.005 ;
        RECT  2.475 2.280 2.755 2.735 ;
        RECT  2.245 1.775 2.610 2.005 ;
        RECT  2.015 1.775 2.245 3.265 ;
        RECT  2.115 1.040 2.170 1.380 ;
        RECT  1.830 3.495 2.170 3.835 ;
        RECT  1.830 1.040 2.115 1.400 ;
        RECT  1.780 1.170 1.830 1.400 ;
        RECT  1.780 3.495 1.830 3.725 ;
        RECT  1.550 1.170 1.780 3.725 ;
        RECT  1.085 1.040 1.315 3.865 ;
    END
END MX4X1

MACRO MX2XL
    CLASS CORE ;
    FOREIGN MX2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 1.125 5.140 3.550 ;
        RECT  4.705 1.125 4.910 1.515 ;
        RECT  4.835 3.195 4.910 3.550 ;
        RECT  4.520 3.210 4.835 3.550 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 4.025 0.710 4.400 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.745 1.840 3.220 ;
        RECT  1.100 2.600 1.460 3.065 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 1.760 4.480 2.155 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.295 -0.400 5.280 0.400 ;
        RECT  3.955 -0.400 4.295 0.575 ;
        RECT  1.315 -0.400 3.955 0.400 ;
        RECT  1.315 1.160 1.325 1.500 ;
        RECT  0.995 -0.400 1.315 1.500 ;
        RECT  0.000 -0.400 0.995 0.400 ;
        RECT  0.985 1.160 0.995 1.500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.300 4.640 5.280 5.440 ;
        RECT  3.960 4.465 4.300 5.440 ;
        RECT  1.285 4.640 3.960 5.440 ;
        RECT  1.230 3.455 1.285 5.440 ;
        RECT  0.945 3.295 1.230 5.440 ;
        RECT  0.900 3.295 0.945 3.795 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.445 2.430 4.500 2.770 ;
        RECT  4.160 2.430 4.445 2.840 ;
        RECT  4.135 2.610 4.160 2.840 ;
        RECT  3.905 2.610 4.135 4.065 ;
        RECT  2.990 3.835 3.905 4.065 ;
        RECT  3.480 1.160 3.560 1.505 ;
        RECT  3.250 1.160 3.480 3.440 ;
        RECT  2.760 1.175 2.990 4.065 ;
        RECT  2.505 1.175 2.760 1.405 ;
        RECT  2.530 3.315 2.760 3.705 ;
        RECT  2.300 1.650 2.530 3.025 ;
        RECT  2.125 1.650 2.300 1.880 ;
        RECT  2.070 2.795 2.300 3.805 ;
        RECT  1.895 1.155 2.125 1.880 ;
        RECT  1.660 3.575 2.070 3.805 ;
        RECT  1.735 2.130 2.060 2.515 ;
        RECT  1.785 1.155 1.895 1.495 ;
        RECT  0.465 2.130 1.735 2.360 ;
        RECT  0.465 1.160 0.520 1.500 ;
        RECT  0.465 3.310 0.520 3.650 ;
        RECT  0.235 1.160 0.465 3.650 ;
        RECT  0.180 1.160 0.235 1.500 ;
        RECT  0.180 3.310 0.235 3.650 ;
    END
END MX2XL

MACRO MX2X4
    CLASS CORE ;
    FOREIGN MX2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX2XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 0.700 5.800 3.350 ;
        RECT  5.220 2.970 5.420 3.350 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 2.940 1.840 3.220 ;
        RECT  0.625 2.845 0.975 3.220 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.860 1.770 1.515 2.150 ;
        RECT  0.800 1.820 0.860 2.150 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.625 2.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.410 -0.400 6.600 0.400 ;
        RECT  6.070 -0.400 6.410 0.950 ;
        RECT  5.030 -0.400 6.070 0.400 ;
        RECT  4.690 -0.400 5.030 0.950 ;
        RECT  1.460 -0.400 4.690 0.400 ;
        RECT  1.120 -0.400 1.460 1.540 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.400 4.640 6.600 5.440 ;
        RECT  6.060 4.465 6.400 5.440 ;
        RECT  4.840 4.640 6.060 5.440 ;
        RECT  4.500 4.080 4.840 5.440 ;
        RECT  1.300 4.640 4.500 5.440 ;
        RECT  0.960 3.530 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.340 2.080 6.395 2.420 ;
        RECT  6.110 2.080 6.340 3.840 ;
        RECT  6.055 2.080 6.110 2.420 ;
        RECT  3.370 3.610 6.110 3.840 ;
        RECT  4.855 1.315 5.085 2.735 ;
        RECT  4.060 1.315 4.855 1.545 ;
        RECT  4.010 2.505 4.855 2.735 ;
        RECT  3.780 2.505 4.010 3.310 ;
        RECT  3.600 0.675 3.830 2.130 ;
        RECT  3.670 2.970 3.780 3.310 ;
        RECT  2.040 0.675 3.600 0.905 ;
        RECT  3.140 1.220 3.370 3.840 ;
        RECT  2.610 3.500 3.140 3.840 ;
        RECT  2.600 1.220 2.830 3.185 ;
        RECT  2.275 1.220 2.600 1.560 ;
        RECT  2.375 2.955 2.600 3.185 ;
        RECT  2.145 2.955 2.375 3.745 ;
        RECT  2.040 1.995 2.355 2.340 ;
        RECT  2.080 3.515 2.145 3.745 ;
        RECT  1.740 3.515 2.080 3.855 ;
        RECT  1.810 0.675 2.040 2.610 ;
        RECT  0.395 2.380 1.810 2.610 ;
        RECT  0.395 1.230 0.540 1.570 ;
        RECT  0.395 3.530 0.540 3.870 ;
        RECT  0.165 1.230 0.395 3.870 ;
    END
END MX2X4

MACRO MX2X2
    CLASS CORE ;
    FOREIGN MX2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX2XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.545 0.815 5.775 4.105 ;
        RECT  5.495 0.815 5.545 1.845 ;
        RECT  5.370 2.940 5.545 4.105 ;
        RECT  5.425 0.815 5.495 1.660 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 2.965 1.765 3.195 ;
        RECT  0.835 2.965 1.120 3.340 ;
        RECT  0.780 3.000 0.835 3.340 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.210 1.435 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.770 1.285 5.065 1.515 ;
        RECT  4.535 1.285 4.770 1.540 ;
        RECT  4.305 1.285 4.535 2.415 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.960 -0.400 5.940 0.400 ;
        RECT  4.620 -0.400 4.960 1.000 ;
        RECT  1.510 -0.400 4.620 0.400 ;
        RECT  1.170 -0.400 1.510 1.305 ;
        RECT  0.000 -0.400 1.170 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 4.640 5.940 5.440 ;
        RECT  4.570 4.465 4.910 5.440 ;
        RECT  1.510 4.640 4.570 5.440 ;
        RECT  1.170 3.675 1.510 5.440 ;
        RECT  0.000 4.640 1.170 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.140 2.035 5.255 2.500 ;
        RECT  4.910 2.035 5.140 4.175 ;
        RECT  3.495 3.945 4.910 4.175 ;
        RECT  3.785 1.170 4.015 3.605 ;
        RECT  3.265 1.120 3.495 4.175 ;
        RECT  3.130 1.120 3.265 1.350 ;
        RECT  2.860 3.510 3.265 3.850 ;
        RECT  2.790 1.010 3.130 1.350 ;
        RECT  2.745 1.665 2.975 3.195 ;
        RECT  2.475 1.665 2.745 1.895 ;
        RECT  2.385 2.965 2.745 3.195 ;
        RECT  2.245 0.800 2.475 1.895 ;
        RECT  2.225 2.185 2.455 2.545 ;
        RECT  2.155 2.965 2.385 3.845 ;
        RECT  2.030 0.800 2.245 1.030 ;
        RECT  1.955 2.185 2.225 2.415 ;
        RECT  1.725 1.555 1.955 2.415 ;
        RECT  0.520 1.555 1.725 1.785 ;
        RECT  0.465 3.605 0.540 3.945 ;
        RECT  0.465 1.460 0.520 1.800 ;
        RECT  0.235 1.460 0.465 3.945 ;
        RECT  0.180 1.460 0.235 1.800 ;
        RECT  0.200 3.605 0.235 3.945 ;
    END
END MX2X2

MACRO MX2X1
    CLASS CORE ;
    FOREIGN MX2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 1.125 5.140 3.975 ;
        RECT  4.715 1.125 4.910 1.590 ;
        RECT  4.520 3.165 4.910 3.975 ;
        RECT  4.705 1.125 4.715 1.515 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 3.965 0.710 4.340 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.890 1.840 3.220 ;
        RECT  1.100 2.665 1.460 3.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 1.820 4.480 2.215 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.295 -0.400 5.280 0.400 ;
        RECT  3.955 -0.400 4.295 0.575 ;
        RECT  1.315 -0.400 3.955 0.400 ;
        RECT  1.315 1.160 1.325 1.500 ;
        RECT  0.995 -0.400 1.315 1.500 ;
        RECT  0.000 -0.400 0.995 0.400 ;
        RECT  0.985 1.160 0.995 1.500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.300 4.640 5.280 5.440 ;
        RECT  3.960 4.465 4.300 5.440 ;
        RECT  1.280 4.640 3.960 5.440 ;
        RECT  0.940 3.515 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.160 2.585 4.500 2.925 ;
        RECT  4.135 2.610 4.160 2.925 ;
        RECT  3.905 2.610 4.135 4.065 ;
        RECT  2.990 3.835 3.905 4.065 ;
        RECT  3.250 1.130 3.480 3.520 ;
        RECT  2.760 1.175 2.990 4.065 ;
        RECT  2.465 1.175 2.760 1.405 ;
        RECT  2.530 3.315 2.760 3.705 ;
        RECT  2.300 1.650 2.530 3.025 ;
        RECT  2.085 1.650 2.300 1.880 ;
        RECT  2.070 2.795 2.300 3.725 ;
        RECT  1.855 1.130 2.085 1.880 ;
        RECT  1.660 3.495 2.070 3.725 ;
        RECT  1.735 2.135 2.060 2.515 ;
        RECT  1.745 1.130 1.855 1.470 ;
        RECT  0.465 2.200 1.735 2.430 ;
        RECT  0.465 1.160 0.520 1.500 ;
        RECT  0.465 3.160 0.520 3.500 ;
        RECT  0.235 1.160 0.465 3.500 ;
        RECT  0.180 1.160 0.235 1.500 ;
        RECT  0.180 3.160 0.235 3.500 ;
    END
END MX2X1

MACRO JKFFSRXL
    CLASS CORE ;
    FOREIGN JKFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.170 2.370 7.730 2.750 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.285 1.715 9.515 2.090 ;
        RECT  9.100 1.715 9.285 1.945 ;
        RECT  8.870 1.285 9.100 1.945 ;
        RECT  8.795 1.285 8.870 1.515 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.850 0.865 18.925 2.635 ;
        RECT  18.695 0.865 18.850 3.580 ;
        RECT  18.040 0.865 18.695 1.095 ;
        RECT  18.620 2.405 18.695 3.580 ;
        RECT  18.010 3.350 18.620 3.580 ;
        RECT  18.010 3.900 18.065 4.240 ;
        RECT  17.700 0.665 18.040 1.095 ;
        RECT  17.780 3.350 18.010 4.240 ;
        RECT  17.725 3.900 17.780 4.240 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.485 2.405 19.585 2.635 ;
        RECT  19.485 1.350 19.540 1.845 ;
        RECT  19.485 2.910 19.540 3.470 ;
        RECT  19.255 1.350 19.485 3.470 ;
        RECT  19.200 1.350 19.255 1.845 ;
        RECT  19.200 2.910 19.255 3.470 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 1.790 2.015 2.610 ;
        RECT  1.765 2.380 1.785 2.610 ;
        RECT  1.535 2.380 1.765 2.635 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.490 1.635 3.950 2.165 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 1.790 1.130 2.200 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.780 -0.400 19.800 0.400 ;
        RECT  18.440 -0.400 18.780 0.575 ;
        RECT  17.360 -0.400 18.440 0.400 ;
        RECT  16.940 -0.400 17.360 0.950 ;
        RECT  14.590 -0.400 16.940 0.400 ;
        RECT  14.170 -0.400 14.590 1.050 ;
        RECT  10.895 -0.400 14.170 0.400 ;
        RECT  10.665 -0.400 10.895 1.295 ;
        RECT  7.030 -0.400 10.665 0.400 ;
        RECT  6.690 -0.400 7.030 0.575 ;
        RECT  4.160 -0.400 6.690 0.400 ;
        RECT  3.820 -0.400 4.160 0.575 ;
        RECT  1.680 -0.400 3.820 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.780 4.640 19.800 5.440 ;
        RECT  18.440 3.810 18.780 5.440 ;
        RECT  17.305 4.640 18.440 5.440 ;
        RECT  15.805 4.465 17.305 5.440 ;
        RECT  5.060 4.640 15.805 5.440 ;
        RECT  3.560 4.465 5.060 5.440 ;
        RECT  1.180 4.640 3.560 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.920 2.150 18.200 2.490 ;
        RECT  17.920 1.380 18.080 1.720 ;
        RECT  17.920 2.780 18.065 3.120 ;
        RECT  17.690 1.380 17.920 3.120 ;
        RECT  17.420 2.890 17.690 3.120 ;
        RECT  17.190 2.890 17.420 4.235 ;
        RECT  15.500 4.005 17.190 4.235 ;
        RECT  16.690 1.200 16.920 3.705 ;
        RECT  15.995 1.200 16.690 1.430 ;
        RECT  16.145 3.475 16.690 3.705 ;
        RECT  16.230 1.750 16.460 3.135 ;
        RECT  15.350 1.750 16.230 1.980 ;
        RECT  15.805 3.365 16.145 3.705 ;
        RECT  15.765 1.085 15.995 1.430 ;
        RECT  15.030 3.475 15.805 3.705 ;
        RECT  14.570 2.670 15.775 2.900 ;
        RECT  15.620 1.085 15.765 1.315 ;
        RECT  15.270 4.005 15.500 4.410 ;
        RECT  15.120 1.290 15.350 2.440 ;
        RECT  5.620 4.180 15.270 4.410 ;
        RECT  13.695 1.290 15.120 1.520 ;
        RECT  14.105 2.210 15.120 2.440 ;
        RECT  14.800 3.475 15.030 3.950 ;
        RECT  13.585 1.750 14.830 1.980 ;
        RECT  14.155 3.720 14.800 3.950 ;
        RECT  14.340 2.670 14.570 3.490 ;
        RECT  13.915 3.260 14.340 3.490 ;
        RECT  13.875 2.210 14.105 3.030 ;
        RECT  13.685 3.260 13.915 3.950 ;
        RECT  13.465 0.630 13.695 1.520 ;
        RECT  6.270 3.720 13.685 3.950 ;
        RECT  13.450 1.750 13.585 2.945 ;
        RECT  11.555 0.630 13.465 0.860 ;
        RECT  13.355 1.750 13.450 3.490 ;
        RECT  13.220 2.715 13.355 3.490 ;
        RECT  8.385 3.260 13.220 3.490 ;
        RECT  12.975 2.120 13.125 2.460 ;
        RECT  12.745 2.120 12.975 3.030 ;
        RECT  12.295 2.120 12.745 2.350 ;
        RECT  10.830 2.795 12.745 3.025 ;
        RECT  12.295 1.160 12.350 1.500 ;
        RECT  12.065 1.160 12.295 2.350 ;
        RECT  12.010 1.160 12.065 1.500 ;
        RECT  9.975 2.265 11.790 2.495 ;
        RECT  11.325 0.630 11.555 1.760 ;
        RECT  10.435 1.530 11.325 1.760 ;
        RECT  10.205 0.675 10.435 1.760 ;
        RECT  7.490 0.675 10.205 0.905 ;
        RECT  9.745 1.195 9.975 2.815 ;
        RECT  9.390 1.195 9.745 1.425 ;
        RECT  8.845 2.585 9.745 2.815 ;
        RECT  8.615 2.280 8.845 2.815 ;
        RECT  8.385 1.135 8.450 1.365 ;
        RECT  8.155 1.135 8.385 3.490 ;
        RECT  8.090 1.135 8.155 1.365 ;
        RECT  7.495 3.145 8.155 3.490 ;
        RECT  7.695 1.700 7.925 2.040 ;
        RECT  5.705 1.715 7.695 1.945 ;
        RECT  6.770 3.145 7.495 3.375 ;
        RECT  7.260 0.675 7.490 1.470 ;
        RECT  6.170 1.240 7.260 1.470 ;
        RECT  6.540 2.260 6.770 3.375 ;
        RECT  6.430 2.260 6.540 2.600 ;
        RECT  6.040 3.420 6.270 3.950 ;
        RECT  5.940 0.725 6.170 1.470 ;
        RECT  5.055 3.420 6.040 3.650 ;
        RECT  5.820 0.725 5.940 0.955 ;
        RECT  5.705 2.890 5.860 3.120 ;
        RECT  5.475 1.200 5.705 3.120 ;
        RECT  5.390 3.945 5.620 4.410 ;
        RECT  2.440 3.945 5.390 4.175 ;
        RECT  5.055 1.540 5.180 1.770 ;
        RECT  4.825 1.540 5.055 3.650 ;
        RECT  4.590 1.000 4.960 1.230 ;
        RECT  0.465 3.420 4.825 3.650 ;
        RECT  4.365 2.270 4.595 2.640 ;
        RECT  4.360 1.000 4.590 1.375 ;
        RECT  2.800 2.895 4.500 3.125 ;
        RECT  2.480 2.410 4.365 2.640 ;
        RECT  2.950 1.145 4.360 1.375 ;
        RECT  2.945 1.145 2.950 1.430 ;
        RECT  2.715 1.090 2.945 1.430 ;
        RECT  2.410 1.310 2.480 3.135 ;
        RECT  2.250 1.310 2.410 3.190 ;
        RECT  1.920 1.310 2.250 1.540 ;
        RECT  2.070 2.850 2.250 3.190 ;
        RECT  1.580 1.200 1.920 1.540 ;
        RECT  0.350 1.190 0.465 1.540 ;
        RECT  0.350 2.760 0.465 3.650 ;
        RECT  0.235 1.190 0.350 3.650 ;
        RECT  0.120 1.190 0.235 3.245 ;
    END
END JKFFSRXL

MACRO JKFFSRX4
    CLASS CORE ;
    FOREIGN JKFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSRXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.170 2.370 7.730 2.750 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.285 1.715 9.515 2.210 ;
        RECT  9.100 1.715 9.285 1.945 ;
        RECT  8.820 1.285 9.100 1.945 ;
        RECT  8.795 1.285 8.820 1.515 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.400 1.820 19.660 3.220 ;
        RECT  19.280 1.385 19.400 3.220 ;
        RECT  19.115 1.385 19.280 3.175 ;
        RECT  19.060 1.385 19.115 1.725 ;
        RECT  19.060 2.835 19.115 3.175 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.830 1.820 20.980 3.220 ;
        RECT  20.680 1.445 20.830 3.220 ;
        RECT  20.600 1.390 20.680 3.220 ;
        RECT  20.340 1.390 20.600 1.730 ;
        RECT  20.395 2.715 20.600 3.080 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.790 2.015 2.330 ;
        RECT  1.785 1.790 1.840 2.635 ;
        RECT  1.535 2.100 1.785 2.635 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.490 1.550 3.950 2.080 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 1.790 1.130 2.200 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.325 -0.400 21.780 0.400 ;
        RECT  20.985 -0.400 21.325 0.960 ;
        RECT  20.040 -0.400 20.985 0.400 ;
        RECT  19.700 -0.400 20.040 0.995 ;
        RECT  18.680 -0.400 19.700 0.400 ;
        RECT  18.340 -0.400 18.680 0.960 ;
        RECT  17.275 -0.400 18.340 0.400 ;
        RECT  16.935 -0.400 17.275 1.355 ;
        RECT  14.470 -0.400 16.935 0.400 ;
        RECT  14.050 -0.400 14.470 0.825 ;
        RECT  10.895 -0.400 14.050 0.400 ;
        RECT  10.665 -0.400 10.895 1.510 ;
        RECT  7.030 -0.400 10.665 0.400 ;
        RECT  6.690 -0.400 7.030 0.575 ;
        RECT  4.260 -0.400 6.690 0.400 ;
        RECT  3.920 -0.400 4.260 0.575 ;
        RECT  1.680 -0.400 3.920 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.320 4.640 21.780 5.440 ;
        RECT  20.980 4.010 21.320 5.440 ;
        RECT  20.040 4.640 20.980 5.440 ;
        RECT  19.700 3.970 20.040 5.440 ;
        RECT  18.680 4.640 19.700 5.440 ;
        RECT  18.340 3.980 18.680 5.440 ;
        RECT  17.305 4.640 18.340 5.440 ;
        RECT  16.025 4.465 17.305 5.440 ;
        RECT  5.060 4.640 16.025 5.440 ;
        RECT  3.560 4.465 5.060 5.440 ;
        RECT  1.180 4.640 3.560 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.120 2.045 20.310 2.385 ;
        RECT  19.970 2.045 20.120 3.680 ;
        RECT  19.890 2.100 19.970 3.680 ;
        RECT  18.140 3.450 19.890 3.680 ;
        RECT  18.085 2.740 18.140 3.680 ;
        RECT  18.085 1.460 18.120 1.800 ;
        RECT  18.030 1.460 18.085 3.680 ;
        RECT  17.855 1.460 18.030 4.235 ;
        RECT  17.780 1.460 17.855 1.800 ;
        RECT  17.800 2.740 17.855 4.235 ;
        RECT  15.500 4.005 17.800 4.235 ;
        RECT  16.730 1.620 16.960 3.660 ;
        RECT  15.860 1.620 16.730 1.850 ;
        RECT  16.220 3.430 16.730 3.660 ;
        RECT  16.270 2.100 16.500 2.850 ;
        RECT  15.395 2.100 16.270 2.330 ;
        RECT  15.880 3.430 16.220 3.770 ;
        RECT  14.985 3.540 15.880 3.770 ;
        RECT  14.515 2.565 15.875 2.795 ;
        RECT  15.630 1.000 15.860 1.850 ;
        RECT  15.500 1.000 15.630 1.340 ;
        RECT  15.270 4.005 15.500 4.410 ;
        RECT  15.230 1.590 15.395 2.330 ;
        RECT  5.620 4.180 15.270 4.410 ;
        RECT  15.000 1.055 15.230 2.335 ;
        RECT  13.520 1.055 15.000 1.285 ;
        RECT  14.055 2.105 15.000 2.335 ;
        RECT  14.755 3.540 14.985 3.830 ;
        RECT  13.585 1.645 14.770 1.875 ;
        RECT  14.510 3.600 14.755 3.830 ;
        RECT  14.285 2.565 14.515 3.370 ;
        RECT  14.280 3.600 14.510 3.950 ;
        RECT  14.050 3.140 14.285 3.370 ;
        RECT  13.825 2.105 14.055 2.910 ;
        RECT  13.820 3.140 14.050 3.950 ;
        RECT  6.140 3.720 13.820 3.950 ;
        RECT  13.355 1.645 13.585 3.490 ;
        RECT  13.290 0.630 13.520 1.285 ;
        RECT  8.385 3.260 13.355 3.490 ;
        RECT  11.355 0.630 13.290 0.860 ;
        RECT  12.895 1.520 13.125 3.030 ;
        RECT  12.270 1.520 12.895 1.750 ;
        RECT  10.720 2.800 12.895 3.030 ;
        RECT  11.930 1.335 12.270 1.750 ;
        RECT  11.630 2.205 11.970 2.545 ;
        RECT  9.975 2.260 11.630 2.525 ;
        RECT  11.125 0.630 11.355 1.985 ;
        RECT  10.435 1.755 11.125 1.985 ;
        RECT  10.205 0.675 10.435 1.985 ;
        RECT  7.490 0.675 10.205 0.905 ;
        RECT  9.745 1.250 9.975 3.030 ;
        RECT  9.730 1.250 9.745 1.480 ;
        RECT  8.845 2.800 9.745 3.030 ;
        RECT  9.390 1.140 9.730 1.480 ;
        RECT  8.615 2.280 8.845 3.030 ;
        RECT  8.385 1.195 8.450 1.425 ;
        RECT  8.155 1.195 8.385 3.490 ;
        RECT  8.090 1.195 8.155 1.425 ;
        RECT  7.780 3.145 8.155 3.430 ;
        RECT  7.695 1.700 7.925 2.040 ;
        RECT  7.440 3.090 7.780 3.430 ;
        RECT  5.705 1.715 7.695 1.945 ;
        RECT  7.260 0.675 7.490 1.470 ;
        RECT  6.770 3.145 7.440 3.375 ;
        RECT  6.170 1.240 7.260 1.470 ;
        RECT  6.540 2.260 6.770 3.375 ;
        RECT  6.430 2.260 6.540 2.600 ;
        RECT  5.940 0.725 6.170 1.470 ;
        RECT  5.910 3.415 6.140 3.950 ;
        RECT  5.820 0.725 5.940 0.955 ;
        RECT  5.055 3.415 5.910 3.645 ;
        RECT  5.705 2.875 5.860 3.105 ;
        RECT  5.475 1.200 5.705 3.105 ;
        RECT  5.390 3.945 5.620 4.410 ;
        RECT  3.380 3.945 5.390 4.175 ;
        RECT  5.055 1.470 5.165 1.810 ;
        RECT  4.825 1.470 5.055 3.645 ;
        RECT  2.950 0.995 4.960 1.225 ;
        RECT  0.520 3.415 4.825 3.645 ;
        RECT  4.365 2.260 4.595 2.610 ;
        RECT  4.160 2.845 4.500 3.185 ;
        RECT  2.480 2.380 4.365 2.610 ;
        RECT  3.425 2.895 4.160 3.125 ;
        RECT  3.195 2.845 3.425 3.125 ;
        RECT  2.440 3.890 3.380 4.230 ;
        RECT  2.760 2.845 3.195 3.075 ;
        RECT  2.945 0.995 2.950 1.280 ;
        RECT  2.715 0.940 2.945 1.280 ;
        RECT  2.250 1.310 2.480 3.175 ;
        RECT  1.920 1.310 2.250 1.540 ;
        RECT  2.060 2.945 2.250 3.175 ;
        RECT  1.580 1.200 1.920 1.540 ;
        RECT  0.410 2.880 0.520 3.645 ;
        RECT  0.350 1.190 0.465 1.540 ;
        RECT  0.350 2.460 0.410 3.645 ;
        RECT  0.290 1.190 0.350 3.645 ;
        RECT  0.180 1.190 0.290 3.220 ;
        RECT  0.120 1.190 0.180 2.690 ;
    END
END JKFFSRX4

MACRO JKFFSRX2
    CLASS CORE ;
    FOREIGN JKFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSRXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.170 2.370 7.730 2.750 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.285 1.715 9.515 2.210 ;
        RECT  9.100 1.715 9.285 1.945 ;
        RECT  8.870 1.285 9.100 1.945 ;
        RECT  8.795 1.285 8.870 1.515 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.765 2.405 18.925 3.080 ;
        RECT  18.765 0.765 18.820 1.575 ;
        RECT  18.535 0.765 18.765 3.080 ;
        RECT  18.480 0.765 18.535 1.575 ;
        RECT  18.500 2.740 18.535 3.080 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.245 2.620 20.280 4.220 ;
        RECT  20.205 0.765 20.260 1.575 ;
        RECT  20.205 2.405 20.245 4.220 ;
        RECT  19.975 0.765 20.205 4.220 ;
        RECT  19.920 0.765 19.975 1.575 ;
        RECT  19.940 2.620 19.975 4.220 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.790 2.015 2.330 ;
        RECT  1.785 1.790 1.840 2.635 ;
        RECT  1.535 2.100 1.785 2.635 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.490 1.550 3.950 2.080 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 1.790 1.130 2.200 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.540 -0.400 20.460 0.400 ;
        RECT  19.200 -0.400 19.540 1.575 ;
        RECT  17.275 -0.400 19.200 0.400 ;
        RECT  16.935 -0.400 17.275 0.575 ;
        RECT  14.470 -0.400 16.935 0.400 ;
        RECT  14.050 -0.400 14.470 0.825 ;
        RECT  10.895 -0.400 14.050 0.400 ;
        RECT  10.665 -0.400 10.895 1.510 ;
        RECT  7.030 -0.400 10.665 0.400 ;
        RECT  6.690 -0.400 7.030 0.575 ;
        RECT  4.260 -0.400 6.690 0.400 ;
        RECT  3.920 -0.400 4.260 0.575 ;
        RECT  1.680 -0.400 3.920 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.560 4.640 20.460 5.440 ;
        RECT  19.220 3.950 19.560 5.440 ;
        RECT  17.305 4.640 19.220 5.440 ;
        RECT  16.025 4.465 17.305 5.440 ;
        RECT  5.060 4.640 16.025 5.440 ;
        RECT  3.560 4.465 5.060 5.440 ;
        RECT  1.180 4.640 3.560 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.465 2.045 19.695 3.680 ;
        RECT  18.140 3.450 19.465 3.680 ;
        RECT  18.085 2.895 18.140 3.705 ;
        RECT  18.085 1.170 18.120 1.510 ;
        RECT  18.030 1.170 18.085 3.705 ;
        RECT  17.855 1.170 18.030 4.235 ;
        RECT  17.780 1.170 17.855 1.510 ;
        RECT  17.800 2.895 17.855 4.235 ;
        RECT  15.500 4.005 17.800 4.235 ;
        RECT  16.800 1.110 17.030 3.775 ;
        RECT  15.840 1.110 16.800 1.340 ;
        RECT  14.985 3.545 16.800 3.775 ;
        RECT  16.445 2.510 16.555 2.850 ;
        RECT  16.215 1.645 16.445 2.850 ;
        RECT  15.230 1.645 16.215 1.875 ;
        RECT  15.535 2.510 15.875 2.850 ;
        RECT  15.500 1.000 15.840 1.340 ;
        RECT  14.515 2.620 15.535 2.850 ;
        RECT  15.270 4.005 15.500 4.410 ;
        RECT  5.620 4.180 15.270 4.410 ;
        RECT  15.000 1.055 15.230 2.335 ;
        RECT  13.520 1.055 15.000 1.285 ;
        RECT  14.055 2.105 15.000 2.335 ;
        RECT  14.755 3.545 14.985 3.830 ;
        RECT  13.585 1.645 14.770 1.875 ;
        RECT  14.510 3.600 14.755 3.830 ;
        RECT  14.285 2.620 14.515 3.370 ;
        RECT  14.280 3.600 14.510 3.950 ;
        RECT  14.050 3.140 14.285 3.370 ;
        RECT  13.825 2.105 14.055 2.910 ;
        RECT  13.820 3.140 14.050 3.950 ;
        RECT  6.140 3.720 13.820 3.950 ;
        RECT  13.355 1.645 13.585 3.490 ;
        RECT  13.290 0.630 13.520 1.285 ;
        RECT  8.385 3.260 13.355 3.490 ;
        RECT  11.355 0.630 13.290 0.860 ;
        RECT  12.895 1.515 13.125 3.030 ;
        RECT  12.270 1.515 12.895 1.745 ;
        RECT  10.720 2.800 12.895 3.030 ;
        RECT  11.930 1.330 12.270 1.745 ;
        RECT  11.630 2.195 11.970 2.535 ;
        RECT  9.975 2.305 11.630 2.535 ;
        RECT  11.125 0.630 11.355 2.065 ;
        RECT  10.435 1.835 11.125 2.065 ;
        RECT  10.205 0.675 10.435 2.065 ;
        RECT  7.490 0.675 10.205 0.905 ;
        RECT  9.745 1.250 9.975 3.030 ;
        RECT  9.730 1.250 9.745 1.480 ;
        RECT  8.845 2.800 9.745 3.030 ;
        RECT  9.390 1.140 9.730 1.480 ;
        RECT  8.615 2.280 8.845 3.030 ;
        RECT  8.155 1.140 8.385 3.490 ;
        RECT  7.440 3.090 8.155 3.430 ;
        RECT  7.695 1.700 7.925 2.040 ;
        RECT  5.705 1.715 7.695 1.945 ;
        RECT  7.260 0.675 7.490 1.470 ;
        RECT  6.770 3.090 7.440 3.320 ;
        RECT  6.170 1.240 7.260 1.470 ;
        RECT  6.540 2.260 6.770 3.320 ;
        RECT  6.430 2.260 6.540 2.600 ;
        RECT  5.940 0.725 6.170 1.470 ;
        RECT  5.910 3.415 6.140 3.950 ;
        RECT  5.820 0.725 5.940 0.955 ;
        RECT  5.055 3.415 5.910 3.645 ;
        RECT  5.705 2.820 5.860 3.160 ;
        RECT  5.475 1.200 5.705 3.160 ;
        RECT  5.390 3.945 5.620 4.410 ;
        RECT  3.380 3.945 5.390 4.175 ;
        RECT  5.055 1.525 5.180 1.755 ;
        RECT  4.825 1.525 5.055 3.645 ;
        RECT  4.840 0.935 4.960 1.165 ;
        RECT  4.610 0.935 4.840 1.225 ;
        RECT  0.520 3.415 4.825 3.645 ;
        RECT  2.950 0.995 4.610 1.225 ;
        RECT  4.365 2.260 4.595 2.610 ;
        RECT  4.160 2.840 4.500 3.180 ;
        RECT  2.480 2.380 4.365 2.610 ;
        RECT  3.375 2.895 4.160 3.125 ;
        RECT  2.440 3.890 3.380 4.230 ;
        RECT  3.145 2.845 3.375 3.125 ;
        RECT  2.760 2.845 3.145 3.075 ;
        RECT  2.945 0.995 2.950 1.280 ;
        RECT  2.715 0.940 2.945 1.280 ;
        RECT  2.250 1.310 2.480 3.175 ;
        RECT  1.920 1.310 2.250 1.540 ;
        RECT  2.060 2.945 2.250 3.175 ;
        RECT  1.580 1.200 1.920 1.540 ;
        RECT  0.350 1.200 0.520 1.540 ;
        RECT  0.350 2.880 0.520 3.645 ;
        RECT  0.290 1.200 0.350 3.645 ;
        RECT  0.120 1.200 0.290 3.220 ;
    END
END JKFFSRX2

MACRO JKFFSRX1
    CLASS CORE ;
    FOREIGN JKFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.170 2.370 7.730 2.750 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.285 1.715 9.515 2.090 ;
        RECT  9.100 1.715 9.285 1.945 ;
        RECT  8.870 1.285 9.100 1.945 ;
        RECT  8.795 1.285 8.870 1.515 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.850 1.845 18.925 2.075 ;
        RECT  18.620 0.865 18.850 3.580 ;
        RECT  18.035 0.865 18.620 1.095 ;
        RECT  18.010 3.350 18.620 3.580 ;
        RECT  17.920 0.725 18.035 1.095 ;
        RECT  17.780 3.350 18.010 4.240 ;
        RECT  17.635 0.665 17.920 1.095 ;
        RECT  17.580 0.665 17.635 1.005 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.485 2.405 19.585 2.635 ;
        RECT  19.255 1.370 19.485 3.600 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 1.790 2.015 2.610 ;
        RECT  1.765 2.380 1.785 2.610 ;
        RECT  1.535 2.380 1.765 2.635 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.490 1.550 3.950 2.080 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 1.790 1.130 2.200 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.780 -0.400 19.800 0.400 ;
        RECT  18.440 -0.400 18.780 0.575 ;
        RECT  17.240 -0.400 18.440 0.400 ;
        RECT  16.820 -0.400 17.240 0.980 ;
        RECT  14.470 -0.400 16.820 0.400 ;
        RECT  14.050 -0.400 14.470 1.060 ;
        RECT  10.895 -0.400 14.050 0.400 ;
        RECT  10.665 -0.400 10.895 1.295 ;
        RECT  7.030 -0.400 10.665 0.400 ;
        RECT  6.690 -0.400 7.030 0.575 ;
        RECT  4.260 -0.400 6.690 0.400 ;
        RECT  3.920 -0.400 4.260 0.575 ;
        RECT  1.680 -0.400 3.920 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.725 4.640 19.800 5.440 ;
        RECT  18.725 3.810 18.780 4.040 ;
        RECT  18.495 3.810 18.725 5.440 ;
        RECT  18.440 3.810 18.495 4.040 ;
        RECT  17.270 4.640 18.495 5.440 ;
        RECT  15.770 4.465 17.270 5.440 ;
        RECT  5.060 4.640 15.770 5.440 ;
        RECT  3.560 4.465 5.060 5.440 ;
        RECT  1.180 4.640 3.560 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.920 2.150 18.200 2.490 ;
        RECT  17.920 2.780 18.065 3.120 ;
        RECT  17.690 1.440 17.920 3.120 ;
        RECT  17.580 1.440 17.690 1.780 ;
        RECT  17.420 2.890 17.690 3.120 ;
        RECT  17.190 2.890 17.420 4.235 ;
        RECT  15.425 4.005 17.190 4.235 ;
        RECT  16.730 1.215 16.960 3.485 ;
        RECT  15.500 1.215 16.730 1.445 ;
        RECT  16.185 3.255 16.730 3.485 ;
        RECT  16.270 1.750 16.500 2.955 ;
        RECT  15.330 1.750 16.270 1.980 ;
        RECT  15.955 3.255 16.185 3.775 ;
        RECT  15.860 3.490 15.955 3.775 ;
        RECT  14.965 3.545 15.860 3.775 ;
        RECT  14.505 2.670 15.785 2.900 ;
        RECT  15.195 4.005 15.425 4.410 ;
        RECT  15.230 1.750 15.330 2.440 ;
        RECT  15.100 1.290 15.230 2.440 ;
        RECT  5.620 4.180 15.195 4.410 ;
        RECT  15.000 1.290 15.100 1.980 ;
        RECT  14.045 2.210 15.100 2.440 ;
        RECT  13.575 1.290 15.000 1.520 ;
        RECT  14.735 3.545 14.965 3.950 ;
        RECT  13.585 1.750 14.770 1.980 ;
        RECT  14.155 3.720 14.735 3.950 ;
        RECT  14.275 2.670 14.505 3.490 ;
        RECT  13.915 3.260 14.275 3.490 ;
        RECT  13.815 2.210 14.045 3.030 ;
        RECT  13.685 3.260 13.915 3.950 ;
        RECT  6.140 3.720 13.685 3.950 ;
        RECT  13.450 1.750 13.585 2.680 ;
        RECT  13.345 0.630 13.575 1.520 ;
        RECT  13.355 1.750 13.450 3.490 ;
        RECT  13.220 2.450 13.355 3.490 ;
        RECT  11.555 0.630 13.345 0.860 ;
        RECT  8.385 3.260 13.220 3.490 ;
        RECT  12.990 1.880 13.125 2.220 ;
        RECT  12.760 1.880 12.990 3.030 ;
        RECT  12.270 1.880 12.760 2.110 ;
        RECT  11.115 2.800 12.760 3.030 ;
        RECT  12.040 1.305 12.270 2.110 ;
        RECT  11.930 1.305 12.040 1.535 ;
        RECT  9.975 2.155 11.790 2.385 ;
        RECT  11.325 0.630 11.555 1.760 ;
        RECT  10.435 1.530 11.325 1.760 ;
        RECT  10.885 2.795 11.115 3.030 ;
        RECT  10.830 2.795 10.885 3.025 ;
        RECT  10.205 0.675 10.435 1.760 ;
        RECT  7.490 0.675 10.205 0.905 ;
        RECT  9.745 1.195 9.975 2.815 ;
        RECT  9.390 1.195 9.745 1.425 ;
        RECT  8.845 2.585 9.745 2.815 ;
        RECT  8.615 2.280 8.845 2.815 ;
        RECT  8.385 1.135 8.450 1.365 ;
        RECT  8.155 1.135 8.385 3.490 ;
        RECT  8.090 1.135 8.155 1.365 ;
        RECT  7.495 3.145 8.155 3.490 ;
        RECT  7.695 1.700 7.925 2.040 ;
        RECT  5.705 1.715 7.695 1.945 ;
        RECT  6.770 3.145 7.495 3.375 ;
        RECT  7.260 0.675 7.490 1.470 ;
        RECT  6.170 1.240 7.260 1.470 ;
        RECT  6.540 2.260 6.770 3.375 ;
        RECT  6.430 2.260 6.540 2.600 ;
        RECT  5.940 0.725 6.170 1.470 ;
        RECT  5.910 3.415 6.140 3.950 ;
        RECT  5.820 0.725 5.940 0.955 ;
        RECT  5.055 3.415 5.910 3.645 ;
        RECT  5.705 2.875 5.860 3.105 ;
        RECT  5.475 1.200 5.705 3.105 ;
        RECT  5.390 3.945 5.620 4.410 ;
        RECT  2.440 3.945 5.390 4.175 ;
        RECT  5.055 1.525 5.180 1.755 ;
        RECT  4.825 1.525 5.055 3.645 ;
        RECT  4.840 0.935 4.960 1.165 ;
        RECT  4.610 0.935 4.840 1.225 ;
        RECT  0.465 3.415 4.825 3.645 ;
        RECT  2.950 0.995 4.610 1.225 ;
        RECT  4.365 2.270 4.595 2.610 ;
        RECT  2.760 2.895 4.500 3.125 ;
        RECT  2.480 2.380 4.365 2.610 ;
        RECT  2.945 0.995 2.950 1.280 ;
        RECT  2.715 0.940 2.945 1.280 ;
        RECT  2.250 1.310 2.480 3.120 ;
        RECT  1.920 1.310 2.250 1.540 ;
        RECT  2.060 2.890 2.250 3.120 ;
        RECT  1.580 1.200 1.920 1.540 ;
        RECT  0.350 1.190 0.465 1.540 ;
        RECT  0.350 2.880 0.465 3.645 ;
        RECT  0.235 1.190 0.350 3.645 ;
        RECT  0.120 1.190 0.235 3.245 ;
    END
END JKFFSRX1

MACRO JKFFSXL
    CLASS CORE ;
    FOREIGN JKFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.900 1.285 12.985 1.515 ;
        RECT  12.670 0.810 12.900 2.040 ;
        RECT  11.990 0.810 12.670 1.040 ;
        RECT  11.760 0.630 11.990 1.040 ;
        RECT  11.665 0.630 11.760 0.980 ;
        RECT  7.475 0.630 11.665 0.860 ;
        RECT  7.425 0.630 7.475 0.955 ;
        RECT  7.195 0.630 7.425 1.700 ;
        RECT  6.860 1.470 7.195 1.700 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.890 2.405 14.965 2.645 ;
        RECT  14.660 1.460 14.890 3.190 ;
        RECT  14.455 1.460 14.660 1.800 ;
        RECT  14.420 2.850 14.660 3.190 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.090 1.460 16.320 3.190 ;
        RECT  15.980 1.460 16.090 1.845 ;
        RECT  15.980 2.405 16.090 3.190 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.725 2.170 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.630 1.755 3.970 2.235 ;
        RECT  3.255 1.755 3.630 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.355 1.105 2.635 ;
        RECT  0.645 1.760 0.875 2.585 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.555 -0.400 16.500 0.400 ;
        RECT  15.215 -0.400 15.555 0.575 ;
        RECT  12.635 -0.400 15.215 0.400 ;
        RECT  12.295 -0.400 12.635 0.575 ;
        RECT  6.945 -0.400 12.295 0.400 ;
        RECT  6.605 -0.400 6.945 1.200 ;
        RECT  4.180 -0.400 6.605 0.400 ;
        RECT  3.840 -0.400 4.180 0.575 ;
        RECT  2.520 -0.400 3.840 0.400 ;
        RECT  2.180 -0.400 2.520 0.575 ;
        RECT  1.120 -0.400 2.180 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.520 4.640 16.500 5.440 ;
        RECT  15.180 4.465 15.520 5.440 ;
        RECT  14.155 4.640 15.180 5.440 ;
        RECT  13.815 4.465 14.155 5.440 ;
        RECT  12.635 4.640 13.815 5.440 ;
        RECT  12.295 4.465 12.635 5.440 ;
        RECT  9.635 4.640 12.295 5.440 ;
        RECT  6.915 4.465 9.635 5.440 ;
        RECT  3.935 4.640 6.915 5.440 ;
        RECT  3.595 4.465 3.935 5.440 ;
        RECT  1.080 4.640 3.595 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.725 0.815 16.110 1.045 ;
        RECT  15.725 3.575 16.110 3.805 ;
        RECT  15.495 0.815 15.725 4.235 ;
        RECT  14.415 0.815 15.495 1.045 ;
        RECT  14.755 4.005 15.495 4.235 ;
        RECT  14.415 3.710 14.755 4.235 ;
        RECT  1.325 4.005 14.415 4.235 ;
        RECT  14.150 2.100 14.320 2.440 ;
        RECT  14.015 2.100 14.150 3.770 ;
        RECT  13.920 1.190 14.015 3.770 ;
        RECT  13.785 1.190 13.920 2.540 ;
        RECT  13.055 3.540 13.920 3.770 ;
        RECT  13.675 1.190 13.785 1.530 ;
        RECT  12.510 2.310 13.785 2.540 ;
        RECT  13.350 2.945 13.690 3.285 ;
        RECT  12.045 3.000 13.350 3.230 ;
        RECT  12.280 2.310 12.510 2.715 ;
        RECT  11.880 2.430 12.045 3.775 ;
        RECT  11.815 1.270 11.880 3.775 ;
        RECT  11.650 1.270 11.815 2.660 ;
        RECT  10.985 3.545 11.815 3.775 ;
        RECT  11.520 1.270 11.650 1.500 ;
        RECT  11.410 2.935 11.575 3.165 ;
        RECT  11.290 1.215 11.520 1.500 ;
        RECT  11.180 1.750 11.410 3.165 ;
        RECT  10.895 1.215 11.290 1.445 ;
        RECT  10.650 1.750 11.180 1.980 ;
        RECT  10.745 2.365 10.905 2.705 ;
        RECT  10.565 2.365 10.745 3.775 ;
        RECT  10.420 1.215 10.650 1.980 ;
        RECT  10.515 2.420 10.565 3.775 ;
        RECT  9.620 2.420 10.515 2.650 ;
        RECT  5.260 3.545 10.515 3.775 ;
        RECT  8.835 1.215 10.420 1.445 ;
        RECT  9.780 2.925 10.235 3.155 ;
        RECT  9.550 2.925 9.780 3.315 ;
        RECT  9.390 2.095 9.620 2.650 ;
        RECT  8.365 3.085 9.550 3.315 ;
        RECT  8.835 2.620 9.135 2.850 ;
        RECT  8.605 1.215 8.835 2.850 ;
        RECT  8.135 1.095 8.365 3.315 ;
        RECT  7.970 1.095 8.135 1.325 ;
        RECT  6.855 2.935 8.135 3.165 ;
        RECT  7.665 1.755 7.895 2.160 ;
        RECT  5.840 1.930 7.665 2.160 ;
        RECT  6.625 2.400 6.855 3.165 ;
        RECT  6.505 2.400 6.625 2.630 ;
        RECT  5.610 0.630 5.840 3.240 ;
        RECT  5.245 0.630 5.610 0.860 ;
        RECT  5.260 1.895 5.315 2.235 ;
        RECT  5.030 1.895 5.260 3.775 ;
        RECT  4.975 1.895 5.030 2.235 ;
        RECT  0.520 3.545 5.030 3.775 ;
        RECT  4.660 0.630 4.885 0.860 ;
        RECT  4.430 0.630 4.660 1.035 ;
        RECT  4.355 1.895 4.585 2.725 ;
        RECT  2.790 2.955 4.535 3.185 ;
        RECT  3.430 0.805 4.430 1.035 ;
        RECT  2.660 2.495 4.355 2.725 ;
        RECT  3.200 0.630 3.430 1.035 ;
        RECT  2.880 0.630 3.200 0.860 ;
        RECT  2.430 1.225 2.660 2.725 ;
        RECT  1.580 1.225 2.430 1.455 ;
        RECT  2.355 2.495 2.430 2.725 ;
        RECT  2.125 2.495 2.355 3.120 ;
        RECT  0.410 1.190 0.520 1.530 ;
        RECT  0.410 2.880 0.520 3.775 ;
        RECT  0.290 1.190 0.410 3.775 ;
        RECT  0.180 1.190 0.290 3.220 ;
    END
END JKFFSXL

MACRO JKFFSX4
    CLASS CORE ;
    FOREIGN JKFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.375 1.285 15.625 1.515 ;
        RECT  15.375 2.120 15.430 2.460 ;
        RECT  15.145 0.810 15.375 2.460 ;
        RECT  12.350 0.810 15.145 1.040 ;
        RECT  15.090 2.120 15.145 2.460 ;
        RECT  12.120 0.630 12.350 1.040 ;
        RECT  11.130 0.630 12.120 0.860 ;
        RECT  10.900 0.630 11.130 1.035 ;
        RECT  9.070 0.805 10.900 1.035 ;
        RECT  8.840 0.735 9.070 1.035 ;
        RECT  6.905 0.735 8.840 0.965 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.300 1.260 18.340 2.660 ;
        RECT  17.880 1.260 18.300 3.065 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.260 1.260 19.680 3.065 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.725 2.170 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.255 1.755 3.970 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 2.225 1.105 2.635 ;
        RECT  0.645 2.040 0.880 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.280 -0.400 20.460 0.400 ;
        RECT  19.940 -0.400 20.280 0.950 ;
        RECT  18.955 -0.400 19.940 0.400 ;
        RECT  18.615 -0.400 18.955 0.950 ;
        RECT  17.610 -0.400 18.615 0.400 ;
        RECT  17.270 -0.400 17.610 0.950 ;
        RECT  15.820 -0.400 17.270 0.400 ;
        RECT  15.480 -0.400 15.820 0.575 ;
        RECT  13.180 -0.400 15.480 0.400 ;
        RECT  12.840 -0.400 13.180 0.575 ;
        RECT  10.145 -0.400 12.840 0.400 ;
        RECT  9.805 -0.400 10.145 0.575 ;
        RECT  6.670 -0.400 9.805 0.400 ;
        RECT  6.330 -0.400 6.670 0.915 ;
        RECT  4.150 -0.400 6.330 0.400 ;
        RECT  3.810 -0.400 4.150 0.575 ;
        RECT  2.490 -0.400 3.810 0.400 ;
        RECT  2.150 -0.400 2.490 0.575 ;
        RECT  1.090 -0.400 2.150 0.400 ;
        RECT  0.750 -0.400 1.090 0.575 ;
        RECT  0.000 -0.400 0.750 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.280 4.640 20.460 5.440 ;
        RECT  19.940 3.860 20.280 5.440 ;
        RECT  18.955 4.640 19.940 5.440 ;
        RECT  18.615 3.860 18.955 5.440 ;
        RECT  17.580 4.640 18.615 5.440 ;
        RECT  17.240 3.860 17.580 5.440 ;
        RECT  16.050 4.640 17.240 5.440 ;
        RECT  15.710 4.465 16.050 5.440 ;
        RECT  13.015 4.640 15.710 5.440 ;
        RECT  12.675 4.465 13.015 5.440 ;
        RECT  9.515 4.640 12.675 5.440 ;
        RECT  6.795 4.465 9.515 5.440 ;
        RECT  3.890 4.640 6.795 5.440 ;
        RECT  3.550 4.465 3.890 5.440 ;
        RECT  1.080 4.640 3.550 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.195 2.210 20.250 2.550 ;
        RECT  19.965 2.210 20.195 3.585 ;
        RECT  19.910 2.210 19.965 2.550 ;
        RECT  17.630 3.355 19.965 3.585 ;
        RECT  17.400 1.420 17.630 3.585 ;
        RECT  16.900 1.420 17.400 1.650 ;
        RECT  16.845 2.750 17.400 3.095 ;
        RECT  16.800 2.020 17.140 2.360 ;
        RECT  16.560 1.310 16.900 1.650 ;
        RECT  16.615 2.750 16.845 4.235 ;
        RECT  16.145 2.075 16.800 2.305 ;
        RECT  16.560 2.750 16.615 3.090 ;
        RECT  1.325 4.005 16.615 4.235 ;
        RECT  15.915 2.075 16.145 3.645 ;
        RECT  14.745 3.415 15.915 3.645 ;
        RECT  14.515 1.825 14.745 3.645 ;
        RECT  14.500 1.825 14.515 2.055 ;
        RECT  13.470 3.415 14.515 3.645 ;
        RECT  14.160 1.360 14.500 2.055 ;
        RECT  13.920 2.335 14.260 2.675 ;
        RECT  12.335 1.825 14.160 2.055 ;
        RECT  12.195 2.390 13.920 2.620 ;
        RECT  12.065 2.390 12.195 3.775 ;
        RECT  11.965 1.325 12.065 3.775 ;
        RECT  11.835 1.325 11.965 2.620 ;
        RECT  11.090 3.545 11.965 3.775 ;
        RECT  11.615 1.325 11.835 1.555 ;
        RECT  11.575 2.955 11.705 3.185 ;
        RECT  11.385 1.090 11.615 1.555 ;
        RECT  11.345 1.790 11.575 3.185 ;
        RECT  11.235 1.790 11.345 2.130 ;
        RECT  11.150 1.790 11.235 2.020 ;
        RECT  10.920 1.265 11.150 2.020 ;
        RECT  8.825 1.265 10.920 1.495 ;
        RECT  10.685 2.260 10.905 2.600 ;
        RECT  10.455 1.730 10.685 3.775 ;
        RECT  9.510 1.730 10.455 1.960 ;
        RECT  5.045 3.545 10.455 3.775 ;
        RECT  9.950 2.260 10.180 3.315 ;
        RECT  8.365 3.085 9.950 3.315 ;
        RECT  9.280 1.730 9.510 2.300 ;
        RECT  8.825 2.625 9.285 2.855 ;
        RECT  8.595 1.265 8.825 2.855 ;
        RECT  8.135 1.325 8.365 3.315 ;
        RECT  7.815 1.325 8.135 1.555 ;
        RECT  6.855 3.055 8.135 3.315 ;
        RECT  7.665 2.020 7.895 2.495 ;
        RECT  5.690 2.020 7.665 2.250 ;
        RECT  6.625 2.485 6.855 3.315 ;
        RECT  6.385 2.485 6.625 2.715 ;
        RECT  5.460 0.630 5.690 3.300 ;
        RECT  5.215 0.630 5.460 0.860 ;
        RECT  5.045 1.755 5.100 2.095 ;
        RECT  4.815 1.755 5.045 3.775 ;
        RECT  4.630 0.630 4.855 0.860 ;
        RECT  4.760 1.755 4.815 2.095 ;
        RECT  0.520 3.545 4.815 3.775 ;
        RECT  4.400 0.630 4.630 1.035 ;
        RECT  4.355 2.375 4.585 2.765 ;
        RECT  2.790 3.055 4.455 3.285 ;
        RECT  3.400 0.805 4.400 1.035 ;
        RECT  2.665 2.375 4.355 2.605 ;
        RECT  3.170 0.630 3.400 1.035 ;
        RECT  2.850 0.630 3.170 0.860 ;
        RECT  2.435 1.225 2.665 2.605 ;
        RECT  1.550 1.225 2.435 1.455 ;
        RECT  2.355 2.375 2.435 2.605 ;
        RECT  2.125 2.375 2.355 3.120 ;
        RECT  0.410 1.180 0.520 1.520 ;
        RECT  0.410 2.830 0.520 3.775 ;
        RECT  0.290 1.180 0.410 3.775 ;
        RECT  0.180 1.180 0.290 3.170 ;
    END
END JKFFSX4

MACRO JKFFSX2
    CLASS CORE ;
    FOREIGN JKFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.670 0.675 14.550 0.905 ;
        RECT  13.325 0.675 13.670 1.040 ;
        RECT  12.125 0.810 13.325 1.040 ;
        RECT  11.895 0.630 12.125 1.040 ;
        RECT  11.660 0.630 11.895 0.980 ;
        RECT  7.475 0.630 11.660 0.860 ;
        RECT  7.380 0.630 7.475 0.980 ;
        RECT  7.150 0.630 7.380 1.700 ;
        RECT  6.860 1.470 7.150 1.700 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.250 1.455 16.360 2.130 ;
        RECT  16.020 1.455 16.250 2.970 ;
        RECT  15.980 2.635 16.020 2.970 ;
        RECT  15.895 2.740 15.980 2.970 ;
        RECT  15.555 2.740 15.895 3.080 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.300 1.460 17.640 1.800 ;
        RECT  16.945 1.570 17.300 1.800 ;
        RECT  16.945 2.740 17.175 3.265 ;
        RECT  16.715 1.570 16.945 3.265 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.725 2.170 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.255 1.755 3.970 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.355 1.105 2.635 ;
        RECT  0.645 1.760 0.875 2.585 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.000 -0.400 17.820 0.400 ;
        RECT  16.660 -0.400 17.000 1.115 ;
        RECT  15.620 -0.400 16.660 0.400 ;
        RECT  15.280 -0.400 15.620 0.575 ;
        RECT  12.695 -0.400 15.280 0.400 ;
        RECT  12.355 -0.400 12.695 0.575 ;
        RECT  6.915 -0.400 12.355 0.400 ;
        RECT  6.575 -0.400 6.915 1.200 ;
        RECT  4.150 -0.400 6.575 0.400 ;
        RECT  3.810 -0.400 4.150 0.575 ;
        RECT  2.490 -0.400 3.810 0.400 ;
        RECT  2.150 -0.400 2.490 0.575 ;
        RECT  1.090 -0.400 2.150 0.400 ;
        RECT  0.750 -0.400 1.090 0.575 ;
        RECT  0.000 -0.400 0.750 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.535 4.640 17.820 5.440 ;
        RECT  16.195 4.020 16.535 5.440 ;
        RECT  14.395 4.640 16.195 5.440 ;
        RECT  14.055 4.465 14.395 5.440 ;
        RECT  9.635 4.640 14.055 5.440 ;
        RECT  6.915 4.465 9.635 5.440 ;
        RECT  3.935 4.640 6.915 5.440 ;
        RECT  3.595 4.465 3.935 5.440 ;
        RECT  1.080 4.640 3.595 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.410 2.135 17.640 3.775 ;
        RECT  17.210 2.135 17.410 2.475 ;
        RECT  15.155 3.545 17.410 3.775 ;
        RECT  15.045 1.365 15.155 3.775 ;
        RECT  14.925 1.365 15.045 4.235 ;
        RECT  14.895 1.365 14.925 1.595 ;
        RECT  14.815 3.410 14.925 4.235 ;
        RECT  14.555 1.255 14.895 1.595 ;
        RECT  1.325 4.005 14.815 4.235 ;
        RECT  14.490 2.290 14.615 2.630 ;
        RECT  14.260 1.825 14.490 3.505 ;
        RECT  14.195 1.825 14.260 2.055 ;
        RECT  13.175 3.275 14.260 3.505 ;
        RECT  13.855 1.360 14.195 2.055 ;
        RECT  13.555 2.315 13.895 2.655 ;
        RECT  12.120 1.825 13.855 2.055 ;
        RECT  12.165 2.425 13.555 2.655 ;
        RECT  11.935 2.425 12.165 3.775 ;
        RECT  11.880 2.425 11.935 2.655 ;
        RECT  10.985 3.545 11.935 3.775 ;
        RECT  11.650 1.270 11.880 2.655 ;
        RECT  11.410 2.955 11.705 3.185 ;
        RECT  11.520 1.270 11.650 1.500 ;
        RECT  11.290 1.215 11.520 1.500 ;
        RECT  11.180 1.750 11.410 3.185 ;
        RECT  10.895 1.215 11.290 1.445 ;
        RECT  10.650 1.750 11.180 1.980 ;
        RECT  10.745 2.365 10.905 2.705 ;
        RECT  10.565 2.365 10.745 3.775 ;
        RECT  10.420 1.215 10.650 1.980 ;
        RECT  10.515 2.420 10.565 3.775 ;
        RECT  9.620 2.420 10.515 2.650 ;
        RECT  5.260 3.545 10.515 3.775 ;
        RECT  8.835 1.215 10.420 1.445 ;
        RECT  9.780 2.925 10.235 3.155 ;
        RECT  9.550 2.925 9.780 3.315 ;
        RECT  9.390 2.095 9.620 2.650 ;
        RECT  8.365 3.085 9.550 3.315 ;
        RECT  8.835 2.620 9.135 2.850 ;
        RECT  8.605 1.215 8.835 2.850 ;
        RECT  8.135 1.175 8.365 3.315 ;
        RECT  7.940 1.175 8.135 1.405 ;
        RECT  6.855 2.935 8.135 3.165 ;
        RECT  7.665 1.755 7.895 2.160 ;
        RECT  5.840 1.930 7.665 2.160 ;
        RECT  6.625 2.400 6.855 3.165 ;
        RECT  6.505 2.400 6.625 2.630 ;
        RECT  5.610 0.630 5.840 3.195 ;
        RECT  5.215 0.630 5.610 0.860 ;
        RECT  5.260 1.755 5.315 2.095 ;
        RECT  5.030 1.755 5.260 3.775 ;
        RECT  4.975 1.755 5.030 2.095 ;
        RECT  0.520 3.545 5.030 3.775 ;
        RECT  4.630 0.630 4.855 0.860 ;
        RECT  4.400 0.630 4.630 1.035 ;
        RECT  4.355 1.990 4.585 2.605 ;
        RECT  2.790 2.955 4.535 3.185 ;
        RECT  3.400 0.805 4.400 1.035 ;
        RECT  2.630 2.375 4.355 2.605 ;
        RECT  3.170 0.630 3.400 1.035 ;
        RECT  2.850 0.630 3.170 0.860 ;
        RECT  2.400 1.225 2.630 2.610 ;
        RECT  1.550 1.225 2.400 1.455 ;
        RECT  2.355 2.375 2.400 2.610 ;
        RECT  2.125 2.375 2.355 3.120 ;
        RECT  0.410 1.180 0.520 1.520 ;
        RECT  0.410 2.830 0.520 3.775 ;
        RECT  0.290 1.180 0.410 3.775 ;
        RECT  0.180 1.180 0.290 3.170 ;
    END
END JKFFSX2

MACRO JKFFSX1
    CLASS CORE ;
    FOREIGN JKFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.900 1.285 12.985 1.515 ;
        RECT  12.670 0.810 12.900 2.040 ;
        RECT  11.990 0.810 12.670 1.040 ;
        RECT  11.760 0.630 11.990 1.040 ;
        RECT  11.665 0.630 11.760 0.980 ;
        RECT  7.475 0.630 11.665 0.860 ;
        RECT  7.425 0.630 7.475 0.955 ;
        RECT  7.195 0.630 7.425 1.700 ;
        RECT  6.860 1.470 7.195 1.700 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.545 1.380 15.655 1.845 ;
        RECT  15.545 2.980 15.655 3.320 ;
        RECT  15.545 2.405 15.625 2.645 ;
        RECT  15.315 1.380 15.545 3.320 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.750 1.370 16.980 3.320 ;
        RECT  16.640 1.370 16.750 1.845 ;
        RECT  16.715 2.405 16.750 2.635 ;
        RECT  16.640 2.980 16.750 3.320 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.725 2.170 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.255 1.755 3.970 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.355 1.105 2.635 ;
        RECT  0.645 1.760 0.875 2.585 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.215 -0.400 17.160 0.400 ;
        RECT  15.875 -0.400 16.215 0.575 ;
        RECT  14.935 -0.400 15.875 0.400 ;
        RECT  14.595 -0.400 14.935 0.575 ;
        RECT  12.635 -0.400 14.595 0.400 ;
        RECT  12.295 -0.400 12.635 0.575 ;
        RECT  6.945 -0.400 12.295 0.400 ;
        RECT  6.605 -0.400 6.945 1.200 ;
        RECT  4.180 -0.400 6.605 0.400 ;
        RECT  3.840 -0.400 4.180 0.575 ;
        RECT  2.520 -0.400 3.840 0.400 ;
        RECT  2.180 -0.400 2.520 0.575 ;
        RECT  0.640 -0.400 2.180 0.400 ;
        RECT  0.300 -0.400 0.640 0.575 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.415 4.640 17.160 5.440 ;
        RECT  16.075 4.465 16.415 5.440 ;
        RECT  15.115 4.640 16.075 5.440 ;
        RECT  14.515 4.465 15.115 5.440 ;
        RECT  14.155 4.640 14.515 5.440 ;
        RECT  13.815 4.465 14.155 5.440 ;
        RECT  12.635 4.640 13.815 5.440 ;
        RECT  12.295 4.465 12.635 5.440 ;
        RECT  9.635 4.640 12.295 5.440 ;
        RECT  6.915 4.465 9.635 5.440 ;
        RECT  3.935 4.640 6.915 5.440 ;
        RECT  3.595 4.465 3.935 5.440 ;
        RECT  1.080 4.640 3.595 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.400 0.805 16.770 1.035 ;
        RECT  16.400 3.890 16.770 4.120 ;
        RECT  16.170 0.805 16.400 4.235 ;
        RECT  14.880 0.805 16.170 1.035 ;
        RECT  14.945 4.005 16.170 4.235 ;
        RECT  14.695 2.255 15.035 2.595 ;
        RECT  14.605 3.640 14.945 4.235 ;
        RECT  14.650 0.805 14.880 1.470 ;
        RECT  14.150 2.310 14.695 2.540 ;
        RECT  1.325 4.005 14.605 4.235 ;
        RECT  13.975 0.795 14.150 3.775 ;
        RECT  13.920 0.740 13.975 3.775 ;
        RECT  13.635 0.740 13.920 1.080 ;
        RECT  12.510 2.310 13.920 2.540 ;
        RECT  13.055 3.545 13.920 3.775 ;
        RECT  13.350 2.945 13.690 3.285 ;
        RECT  12.045 3.000 13.350 3.230 ;
        RECT  12.280 2.310 12.510 2.715 ;
        RECT  11.880 2.430 12.045 3.775 ;
        RECT  11.815 1.270 11.880 3.775 ;
        RECT  11.650 1.270 11.815 2.660 ;
        RECT  10.985 3.545 11.815 3.775 ;
        RECT  11.520 1.270 11.650 1.500 ;
        RECT  11.410 2.955 11.575 3.185 ;
        RECT  11.290 1.215 11.520 1.500 ;
        RECT  11.180 1.750 11.410 3.185 ;
        RECT  10.895 1.215 11.290 1.445 ;
        RECT  10.650 1.750 11.180 1.980 ;
        RECT  10.745 2.365 10.905 2.705 ;
        RECT  10.565 2.365 10.745 3.775 ;
        RECT  10.420 1.215 10.650 1.980 ;
        RECT  10.515 2.420 10.565 3.775 ;
        RECT  9.620 2.420 10.515 2.650 ;
        RECT  5.260 3.545 10.515 3.775 ;
        RECT  8.835 1.215 10.420 1.445 ;
        RECT  9.780 2.925 10.235 3.155 ;
        RECT  9.550 2.925 9.780 3.315 ;
        RECT  9.390 2.095 9.620 2.650 ;
        RECT  8.365 3.085 9.550 3.315 ;
        RECT  8.835 2.620 9.135 2.850 ;
        RECT  8.605 1.215 8.835 2.850 ;
        RECT  8.135 1.175 8.365 3.315 ;
        RECT  7.970 1.175 8.135 1.405 ;
        RECT  6.855 2.935 8.135 3.165 ;
        RECT  7.665 1.755 7.895 2.160 ;
        RECT  5.840 1.930 7.665 2.160 ;
        RECT  6.625 2.400 6.855 3.165 ;
        RECT  6.505 2.400 6.625 2.630 ;
        RECT  5.610 0.630 5.840 3.195 ;
        RECT  5.245 0.630 5.610 0.860 ;
        RECT  5.260 1.755 5.315 2.095 ;
        RECT  5.030 1.755 5.260 3.775 ;
        RECT  4.975 1.755 5.030 2.095 ;
        RECT  0.520 3.545 5.030 3.775 ;
        RECT  4.660 0.630 4.885 0.860 ;
        RECT  4.430 0.630 4.660 1.035 ;
        RECT  4.355 1.990 4.585 2.605 ;
        RECT  2.790 2.955 4.535 3.185 ;
        RECT  3.430 0.805 4.430 1.035 ;
        RECT  2.660 2.375 4.355 2.605 ;
        RECT  3.200 0.630 3.430 1.035 ;
        RECT  2.880 0.630 3.200 0.860 ;
        RECT  2.630 1.225 2.660 2.605 ;
        RECT  2.430 1.225 2.630 2.610 ;
        RECT  1.580 1.225 2.430 1.455 ;
        RECT  2.355 2.375 2.430 2.610 ;
        RECT  2.125 2.375 2.355 3.120 ;
        RECT  0.410 1.180 0.520 1.520 ;
        RECT  0.410 2.830 0.520 3.775 ;
        RECT  0.290 1.180 0.410 3.775 ;
        RECT  0.180 1.180 0.290 3.170 ;
    END
END JKFFSX1

MACRO JKFFRXL
    CLASS CORE ;
    FOREIGN JKFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.645 1.795 9.100 2.290 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.705 0.770 15.835 1.000 ;
        RECT  15.475 0.770 15.705 1.120 ;
        RECT  15.320 0.890 15.475 1.120 ;
        RECT  15.090 0.890 15.320 3.350 ;
        RECT  14.660 1.260 15.090 1.540 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.745 2.940 17.020 3.220 ;
        RECT  16.645 1.395 16.745 3.320 ;
        RECT  16.515 1.090 16.645 3.320 ;
        RECT  16.360 1.090 16.515 1.715 ;
        RECT  16.355 2.980 16.515 3.320 ;
        RECT  16.305 1.090 16.360 1.430 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.820 1.980 2.405 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 1.935 3.865 2.165 ;
        RECT  3.670 1.260 3.820 1.540 ;
        RECT  3.440 1.260 3.670 2.165 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.015 2.380 1.180 2.660 ;
        RECT  0.880 2.210 1.015 2.660 ;
        RECT  0.785 2.080 0.880 2.660 ;
        RECT  0.645 2.080 0.785 2.440 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.645 -0.400 17.160 0.400 ;
        RECT  16.305 -0.400 16.645 0.575 ;
        RECT  14.775 -0.400 16.305 0.400 ;
        RECT  14.435 -0.400 14.775 0.575 ;
        RECT  13.155 -0.400 14.435 0.400 ;
        RECT  12.815 -0.400 13.155 0.575 ;
        RECT  8.560 -0.400 12.815 0.400 ;
        RECT  8.220 -0.400 8.560 0.980 ;
        RECT  6.960 -0.400 8.220 0.400 ;
        RECT  6.620 -0.400 6.960 1.210 ;
        RECT  2.720 -0.400 6.620 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  1.120 -0.400 2.380 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.135 4.640 17.160 5.440 ;
        RECT  15.795 4.465 16.135 5.440 ;
        RECT  13.345 4.640 15.795 5.440 ;
        RECT  13.005 4.465 13.345 5.440 ;
        RECT  10.615 4.640 13.005 5.440 ;
        RECT  6.695 4.465 10.615 5.440 ;
        RECT  1.765 4.640 6.695 5.440 ;
        RECT  0.945 4.465 1.765 5.440 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.280 2.160 16.285 2.500 ;
        RECT  15.780 2.135 16.280 2.525 ;
        RECT  15.550 1.455 15.780 3.995 ;
        RECT  15.320 3.765 15.550 3.995 ;
        RECT  15.090 3.765 15.320 4.295 ;
        RECT  13.820 4.065 15.090 4.295 ;
        RECT  14.675 2.175 14.825 2.595 ;
        RECT  14.445 1.815 14.675 3.755 ;
        RECT  14.075 1.815 14.445 2.045 ;
        RECT  14.280 3.525 14.445 3.755 ;
        RECT  13.870 2.840 14.210 3.180 ;
        RECT  13.845 1.140 14.075 2.045 ;
        RECT  12.860 2.895 13.870 3.125 ;
        RECT  13.025 1.815 13.845 2.045 ;
        RECT  13.615 0.630 13.820 0.860 ;
        RECT  13.590 4.005 13.820 4.295 ;
        RECT  13.385 0.630 13.615 1.035 ;
        RECT  6.455 4.005 13.590 4.235 ;
        RECT  12.585 0.805 13.385 1.035 ;
        RECT  12.795 1.670 13.025 2.045 ;
        RECT  12.630 2.325 12.860 3.655 ;
        RECT  12.480 2.325 12.630 2.555 ;
        RECT  11.745 3.425 12.630 3.655 ;
        RECT  12.355 0.630 12.585 1.035 ;
        RECT  12.250 1.265 12.480 2.555 ;
        RECT  9.305 0.630 12.355 0.860 ;
        RECT  12.020 2.855 12.275 3.085 ;
        RECT  12.125 1.265 12.250 1.495 ;
        RECT  11.895 1.135 12.125 1.495 ;
        RECT  11.790 1.780 12.020 3.085 ;
        RECT  11.750 1.135 11.895 1.365 ;
        RECT  11.665 1.780 11.790 2.010 ;
        RECT  11.435 1.630 11.665 2.010 ;
        RECT  11.270 2.305 11.500 3.775 ;
        RECT  11.315 1.630 11.435 1.860 ;
        RECT  11.085 1.425 11.315 1.860 ;
        RECT  5.985 3.545 11.270 3.775 ;
        RECT  10.175 1.425 11.085 1.655 ;
        RECT  10.735 2.810 10.845 3.150 ;
        RECT  10.505 2.810 10.735 3.310 ;
        RECT  7.285 3.080 10.505 3.310 ;
        RECT  9.815 1.090 10.175 1.655 ;
        RECT  9.770 2.615 9.870 2.845 ;
        RECT  9.770 1.425 9.815 1.655 ;
        RECT  9.540 1.425 9.770 2.845 ;
        RECT  9.505 2.095 9.540 2.845 ;
        RECT  9.075 0.630 9.305 1.525 ;
        RECT  8.300 2.620 9.165 2.850 ;
        RECT  8.300 1.295 9.075 1.525 ;
        RECT  8.070 1.295 8.300 2.850 ;
        RECT  7.915 1.775 8.070 2.005 ;
        RECT  7.600 1.010 7.760 1.350 ;
        RECT  7.370 1.010 7.600 2.555 ;
        RECT  7.285 2.325 7.370 2.555 ;
        RECT  6.945 2.325 7.285 3.310 ;
        RECT  5.545 1.600 7.120 1.830 ;
        RECT  6.550 2.325 6.945 2.555 ;
        RECT  6.210 2.270 6.550 2.610 ;
        RECT  6.225 4.005 6.455 4.410 ;
        RECT  2.225 4.180 6.225 4.410 ;
        RECT  5.755 3.545 5.985 3.950 ;
        RECT  5.550 3.715 5.755 3.950 ;
        RECT  4.820 3.715 5.550 3.945 ;
        RECT  5.380 0.990 5.545 2.390 ;
        RECT  5.315 0.990 5.380 3.470 ;
        RECT  5.150 2.160 5.315 3.470 ;
        RECT  4.820 1.560 4.980 1.915 ;
        RECT  4.595 0.755 4.825 1.330 ;
        RECT  4.750 1.560 4.820 3.945 ;
        RECT  4.590 1.685 4.750 3.945 ;
        RECT  3.200 0.755 4.595 0.985 ;
        RECT  0.465 3.255 4.590 3.485 ;
        RECT  2.440 2.790 4.355 3.020 ;
        RECT  2.455 3.720 4.115 3.950 ;
        RECT  2.970 0.755 3.200 1.560 ;
        RECT  2.900 1.330 2.970 1.560 ;
        RECT  2.670 1.330 2.900 1.675 ;
        RECT  2.210 1.295 2.440 3.020 ;
        RECT  1.995 3.855 2.225 4.410 ;
        RECT  1.920 1.295 2.210 1.525 ;
        RECT  2.115 2.790 2.210 3.020 ;
        RECT  1.845 3.855 1.995 4.085 ;
        RECT  1.690 0.740 1.920 1.525 ;
        RECT  1.580 0.740 1.690 1.080 ;
        RECT  0.395 1.070 0.520 1.410 ;
        RECT  0.395 2.730 0.465 3.485 ;
        RECT  0.235 1.070 0.395 3.485 ;
        RECT  0.165 1.070 0.235 2.960 ;
    END
END JKFFRXL

MACRO JKFFRX4
    CLASS CORE ;
    FOREIGN JKFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.985 9.380 2.215 ;
        RECT  8.720 1.820 9.100 2.215 ;
        RECT  8.540 1.985 8.720 2.215 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.320 1.460 20.520 1.690 ;
        RECT  20.320 2.830 20.510 3.170 ;
        RECT  20.015 1.460 20.320 3.220 ;
        RECT  19.940 1.820 20.015 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.685 1.405 21.800 1.745 ;
        RECT  21.685 2.830 21.790 3.170 ;
        RECT  21.640 1.405 21.685 3.170 ;
        RECT  21.460 1.405 21.640 3.220 ;
        RECT  21.455 1.460 21.460 3.220 ;
        RECT  21.260 1.820 21.455 3.220 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.625 1.980 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 1.820 3.970 2.250 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.020 2.380 1.180 2.660 ;
        RECT  0.625 2.040 1.020 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.440 -0.400 23.100 0.400 ;
        RECT  22.100 -0.400 22.440 1.015 ;
        RECT  21.160 -0.400 22.100 0.400 ;
        RECT  20.820 -0.400 21.160 1.015 ;
        RECT  19.870 -0.400 20.820 0.400 ;
        RECT  19.530 -0.400 19.870 1.015 ;
        RECT  17.725 -0.400 19.530 0.400 ;
        RECT  17.385 -0.400 17.725 1.230 ;
        RECT  16.280 -0.400 17.385 0.400 ;
        RECT  15.940 -0.400 16.280 0.950 ;
        RECT  14.280 -0.400 15.940 0.400 ;
        RECT  13.940 -0.400 14.280 0.575 ;
        RECT  11.620 -0.400 13.940 0.400 ;
        RECT  11.390 -0.400 11.620 1.280 ;
        RECT  8.575 -0.400 11.390 0.400 ;
        RECT  8.345 -0.400 8.575 0.880 ;
        RECT  7.140 -0.400 8.345 0.400 ;
        RECT  6.800 -0.400 7.140 1.285 ;
        RECT  2.690 -0.400 6.800 0.400 ;
        RECT  2.350 -0.400 2.690 0.575 ;
        RECT  1.080 -0.400 2.350 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.430 4.640 23.100 5.440 ;
        RECT  22.090 4.010 22.430 5.440 ;
        RECT  21.150 4.640 22.090 5.440 ;
        RECT  20.810 4.010 21.150 5.440 ;
        RECT  19.870 4.640 20.810 5.440 ;
        RECT  19.530 4.010 19.870 5.440 ;
        RECT  18.450 4.640 19.530 5.440 ;
        RECT  18.110 4.465 18.450 5.440 ;
        RECT  15.770 4.640 18.110 5.440 ;
        RECT  15.430 4.465 15.770 5.440 ;
        RECT  13.765 4.640 15.430 5.440 ;
        RECT  13.425 4.465 13.765 5.440 ;
        RECT  7.625 4.640 13.425 5.440 ;
        RECT  6.685 4.465 7.625 5.440 ;
        RECT  1.730 4.640 6.685 5.440 ;
        RECT  0.910 4.465 1.730 5.440 ;
        RECT  0.000 4.640 0.910 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.020 2.025 22.250 3.680 ;
        RECT  19.625 3.450 22.020 3.680 ;
        RECT  19.395 1.425 19.625 3.680 ;
        RECT  19.205 1.425 19.395 1.655 ;
        RECT  19.090 3.000 19.395 3.680 ;
        RECT  18.975 1.025 19.205 1.655 ;
        RECT  18.550 1.970 19.160 2.310 ;
        RECT  18.860 3.000 19.090 4.195 ;
        RECT  18.450 1.025 18.975 1.255 ;
        RECT  12.940 3.965 18.860 4.195 ;
        RECT  18.320 1.545 18.550 3.575 ;
        RECT  18.165 0.890 18.450 1.255 ;
        RECT  17.000 1.545 18.320 1.775 ;
        RECT  17.100 3.345 18.320 3.575 ;
        RECT  18.110 0.890 18.165 1.230 ;
        RECT  17.725 2.065 17.955 2.750 ;
        RECT  16.310 2.065 17.725 2.295 ;
        RECT  16.760 3.290 17.100 3.630 ;
        RECT  16.660 0.955 17.000 1.775 ;
        RECT  16.850 2.540 16.970 2.770 ;
        RECT  16.620 2.540 16.850 2.975 ;
        RECT  15.685 1.195 16.660 1.425 ;
        RECT  15.210 2.745 16.620 2.975 ;
        RECT  16.080 2.065 16.310 2.335 ;
        RECT  15.955 2.105 16.080 2.335 ;
        RECT  15.455 0.740 15.685 1.425 ;
        RECT  14.980 1.415 15.210 3.655 ;
        RECT  12.975 1.415 14.980 1.645 ;
        RECT  12.385 3.425 14.980 3.655 ;
        RECT  14.640 2.830 14.750 3.170 ;
        RECT  14.410 2.115 14.640 3.170 ;
        RECT  14.385 0.880 14.635 1.110 ;
        RECT  10.700 2.115 14.410 2.345 ;
        RECT  14.155 0.810 14.385 1.110 ;
        RECT  13.545 0.810 14.155 1.040 ;
        RECT  13.885 2.835 14.075 3.065 ;
        RECT  13.655 2.835 13.885 3.135 ;
        RECT  11.910 2.905 13.655 3.135 ;
        RECT  13.315 0.645 13.545 1.040 ;
        RECT  12.215 0.645 13.315 0.875 ;
        RECT  12.745 1.125 12.975 1.645 ;
        RECT  12.710 3.965 12.940 4.410 ;
        RECT  12.620 1.125 12.745 1.355 ;
        RECT  8.090 4.180 12.710 4.410 ;
        RECT  12.155 3.425 12.385 3.790 ;
        RECT  11.985 0.645 12.215 1.755 ;
        RECT  11.160 1.525 11.985 1.755 ;
        RECT  11.680 2.905 11.910 3.950 ;
        RECT  8.555 3.720 11.680 3.950 ;
        RECT  11.180 2.780 11.410 3.490 ;
        RECT  9.020 3.260 11.180 3.490 ;
        RECT  10.930 0.685 11.160 1.755 ;
        RECT  9.390 0.685 10.930 0.915 ;
        RECT  10.470 1.150 10.700 2.345 ;
        RECT  10.300 1.205 10.470 2.060 ;
        RECT  10.005 1.720 10.300 2.060 ;
        RECT  9.960 1.720 10.005 2.930 ;
        RECT  9.775 1.775 9.960 2.930 ;
        RECT  9.160 0.685 9.390 1.490 ;
        RECT  8.150 2.615 9.200 2.845 ;
        RECT  9.050 1.150 9.160 1.490 ;
        RECT  8.360 1.260 9.050 1.490 ;
        RECT  8.790 3.075 9.020 3.490 ;
        RECT  7.280 3.075 8.790 3.305 ;
        RECT  8.325 3.540 8.555 3.950 ;
        RECT  8.150 1.260 8.360 1.695 ;
        RECT  5.955 3.540 8.325 3.770 ;
        RECT  8.130 1.260 8.150 2.845 ;
        RECT  7.920 1.465 8.130 2.845 ;
        RECT  7.860 4.005 8.090 4.410 ;
        RECT  7.690 1.000 7.865 1.230 ;
        RECT  6.425 4.005 7.860 4.235 ;
        RECT  7.460 1.000 7.690 2.635 ;
        RECT  7.280 2.405 7.460 2.635 ;
        RECT  6.940 2.405 7.280 3.305 ;
        RECT  7.000 1.515 7.230 1.890 ;
        RECT  5.775 1.515 7.000 1.745 ;
        RECT  6.400 2.405 6.940 2.635 ;
        RECT  6.195 4.005 6.425 4.410 ;
        RECT  6.115 2.270 6.400 2.635 ;
        RECT  2.200 4.180 6.195 4.410 ;
        RECT  6.060 2.270 6.115 2.610 ;
        RECT  5.725 3.540 5.955 3.950 ;
        RECT  5.720 1.070 5.775 1.745 ;
        RECT  4.810 3.720 5.725 3.950 ;
        RECT  5.490 1.070 5.720 2.405 ;
        RECT  5.435 1.070 5.490 1.410 ;
        RECT  5.365 2.175 5.490 2.405 ;
        RECT  5.135 2.175 5.365 3.475 ;
        RECT  4.840 1.560 5.070 1.940 ;
        RECT  4.690 0.810 4.920 1.300 ;
        RECT  4.810 1.710 4.840 1.940 ;
        RECT  4.580 1.710 4.810 3.950 ;
        RECT  3.015 0.810 4.690 1.040 ;
        RECT  2.910 3.135 4.580 3.365 ;
        RECT  4.120 2.560 4.350 2.905 ;
        RECT  2.440 2.675 4.120 2.905 ;
        RECT  3.955 3.600 4.095 3.830 ;
        RECT  3.725 3.600 3.955 3.950 ;
        RECT  2.430 3.720 3.725 3.950 ;
        RECT  2.785 0.810 3.015 1.755 ;
        RECT  2.680 3.135 2.910 3.490 ;
        RECT  2.675 1.415 2.785 1.755 ;
        RECT  0.520 3.260 2.680 3.490 ;
        RECT  2.210 0.830 2.440 3.025 ;
        RECT  1.885 0.830 2.210 1.060 ;
        RECT  2.065 2.675 2.210 3.025 ;
        RECT  1.970 3.930 2.200 4.410 ;
        RECT  1.275 3.930 1.970 4.160 ;
        RECT  1.545 0.720 1.885 1.060 ;
        RECT  0.395 1.300 0.520 1.640 ;
        RECT  0.395 2.960 0.520 3.490 ;
        RECT  0.290 1.300 0.395 3.490 ;
        RECT  0.165 1.300 0.290 3.325 ;
    END
END JKFFRX4

MACRO JKFFRX2
    CLASS CORE ;
    FOREIGN JKFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFRXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 1.800 9.760 2.140 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.910 1.820 17.020 2.100 ;
        RECT  16.910 2.635 16.965 3.080 ;
        RECT  16.680 1.335 16.910 3.080 ;
        RECT  16.640 1.820 16.680 2.100 ;
        RECT  16.640 2.635 16.680 3.080 ;
        RECT  16.625 2.740 16.640 3.080 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.280 1.260 18.340 1.540 ;
        RECT  18.245 1.260 18.280 3.025 ;
        RECT  18.050 1.260 18.245 3.080 ;
        RECT  18.035 1.260 18.050 1.845 ;
        RECT  17.905 2.740 18.050 3.080 ;
        RECT  17.960 1.260 18.035 1.680 ;
        RECT  17.905 1.340 17.960 1.680 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.760 2.165 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.875 1.685 4.215 2.045 ;
        RECT  3.820 1.815 3.875 2.045 ;
        RECT  3.515 1.815 3.820 2.100 ;
        RECT  3.440 1.820 3.515 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 2.380 1.180 2.660 ;
        RECT  0.800 1.810 0.910 2.660 ;
        RECT  0.680 1.810 0.800 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 -0.400 18.480 0.400 ;
        RECT  17.265 -0.400 17.605 0.995 ;
        RECT  15.655 -0.400 17.265 0.400 ;
        RECT  15.315 -0.400 15.655 0.575 ;
        RECT  13.685 -0.400 15.315 0.400 ;
        RECT  13.345 -0.400 13.685 0.575 ;
        RECT  8.965 -0.400 13.345 0.400 ;
        RECT  8.625 -0.400 8.965 1.065 ;
        RECT  7.360 -0.400 8.625 0.400 ;
        RECT  7.020 -0.400 7.360 1.235 ;
        RECT  2.720 -0.400 7.020 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  0.640 -0.400 2.380 0.400 ;
        RECT  0.300 -0.400 0.640 0.575 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 4.640 18.480 5.440 ;
        RECT  17.265 4.050 17.605 5.440 ;
        RECT  15.785 4.640 17.265 5.440 ;
        RECT  15.430 4.465 15.785 5.440 ;
        RECT  13.755 4.640 15.430 5.440 ;
        RECT  13.415 4.465 13.755 5.440 ;
        RECT  8.655 4.640 13.415 5.440 ;
        RECT  7.335 4.465 8.655 5.440 ;
        RECT  4.075 4.640 7.335 5.440 ;
        RECT  3.735 4.465 4.075 5.440 ;
        RECT  1.025 4.640 3.735 5.440 ;
        RECT  0.795 3.815 1.025 5.440 ;
        RECT  0.000 4.640 0.795 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.670 2.050 17.820 2.500 ;
        RECT  17.590 2.050 17.670 3.765 ;
        RECT  17.440 2.270 17.590 3.765 ;
        RECT  16.280 3.535 17.440 3.765 ;
        RECT  16.160 1.360 16.280 4.175 ;
        RECT  16.050 1.205 16.160 4.175 ;
        RECT  15.930 1.205 16.050 1.590 ;
        RECT  13.085 3.945 16.050 4.175 ;
        RECT  15.530 2.420 15.815 2.775 ;
        RECT  15.300 0.970 15.530 3.615 ;
        RECT  14.555 0.970 15.300 1.200 ;
        RECT  13.925 3.385 15.300 3.615 ;
        RECT  14.385 2.425 15.065 2.655 ;
        RECT  14.155 1.445 14.385 2.655 ;
        RECT  14.195 0.630 14.320 0.860 ;
        RECT  13.965 0.630 14.195 1.035 ;
        RECT  13.030 1.445 14.155 1.675 ;
        RECT  13.075 0.805 13.965 1.035 ;
        RECT  13.695 1.905 13.925 3.615 ;
        RECT  13.265 1.905 13.695 2.135 ;
        RECT  13.235 2.420 13.465 3.710 ;
        RECT  13.030 2.420 13.235 2.650 ;
        RECT  12.600 3.480 13.235 3.710 ;
        RECT  12.855 3.945 13.085 4.410 ;
        RECT  12.845 0.630 13.075 1.035 ;
        RECT  12.800 1.265 13.030 2.650 ;
        RECT  12.560 2.880 13.000 3.110 ;
        RECT  9.115 4.180 12.855 4.410 ;
        RECT  9.710 0.630 12.845 0.860 ;
        RECT  12.555 1.265 12.800 1.495 ;
        RECT  12.370 3.480 12.600 3.865 ;
        RECT  12.330 1.725 12.560 3.110 ;
        RECT  12.185 1.150 12.555 1.495 ;
        RECT  12.255 3.635 12.370 3.865 ;
        RECT  10.620 1.725 12.330 1.955 ;
        RECT  11.995 2.335 12.100 2.725 ;
        RECT  11.765 2.335 11.995 3.950 ;
        RECT  9.575 3.720 11.765 3.950 ;
        RECT  11.110 2.610 11.340 3.490 ;
        RECT  10.040 3.260 11.110 3.490 ;
        RECT  10.585 2.795 10.705 3.025 ;
        RECT  10.585 1.095 10.620 1.955 ;
        RECT  10.355 1.095 10.585 3.025 ;
        RECT  10.260 1.095 10.355 1.980 ;
        RECT  10.000 1.585 10.260 1.980 ;
        RECT  9.810 3.075 10.040 3.490 ;
        RECT  8.630 2.615 9.885 2.845 ;
        RECT  7.945 3.075 9.810 3.305 ;
        RECT  9.480 0.630 9.710 1.525 ;
        RECT  9.345 3.540 9.575 3.950 ;
        RECT  8.630 1.295 9.480 1.525 ;
        RECT  6.605 3.540 9.345 3.770 ;
        RECT  8.885 4.005 9.115 4.410 ;
        RECT  7.095 4.005 8.885 4.235 ;
        RECT  8.400 1.295 8.630 2.845 ;
        RECT  8.290 1.735 8.400 2.075 ;
        RECT  8.055 1.000 8.165 1.340 ;
        RECT  7.945 1.000 8.055 2.495 ;
        RECT  7.825 1.000 7.945 3.305 ;
        RECT  7.660 2.265 7.825 3.305 ;
        RECT  6.740 2.265 7.660 2.495 ;
        RECT  6.080 1.595 7.510 1.825 ;
        RECT  6.865 4.005 7.095 4.410 ;
        RECT  4.785 4.180 6.865 4.410 ;
        RECT  6.375 3.540 6.605 3.950 ;
        RECT  5.380 3.720 6.375 3.950 ;
        RECT  5.850 1.010 6.080 3.470 ;
        RECT  5.655 1.010 5.850 1.350 ;
        RECT  5.150 1.555 5.380 3.950 ;
        RECT  5.050 1.015 5.190 1.245 ;
        RECT  5.055 1.555 5.150 1.900 ;
        RECT  2.805 2.835 5.150 3.065 ;
        RECT  5.000 1.560 5.055 1.900 ;
        RECT  4.820 0.755 5.050 1.245 ;
        RECT  2.625 2.335 4.920 2.565 ;
        RECT  3.220 0.755 4.820 0.985 ;
        RECT  4.555 3.875 4.785 4.410 ;
        RECT  3.035 3.310 4.775 3.540 ;
        RECT  1.280 3.875 4.555 4.105 ;
        RECT  2.990 0.755 3.220 1.380 ;
        RECT  2.880 1.040 2.990 1.380 ;
        RECT  2.575 2.835 2.805 3.560 ;
        RECT  2.395 1.250 2.625 2.565 ;
        RECT  0.465 3.330 2.575 3.560 ;
        RECT  1.920 1.250 2.395 1.480 ;
        RECT  2.345 2.335 2.395 2.565 ;
        RECT  2.115 2.335 2.345 3.100 ;
        RECT  1.580 1.140 1.920 1.480 ;
        RECT  0.440 1.130 0.520 1.470 ;
        RECT  0.440 2.940 0.465 3.560 ;
        RECT  0.210 1.130 0.440 3.560 ;
        RECT  0.180 1.130 0.210 1.470 ;
    END
END JKFFRX2

MACRO JKFFRX1
    CLASS CORE ;
    FOREIGN JKFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFRXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 1.800 9.760 2.140 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.615 0.735 17.010 1.095 ;
        RECT  16.430 0.865 16.615 1.095 ;
        RECT  16.200 0.865 16.430 3.560 ;
        RECT  15.980 1.820 16.200 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.760 1.350 18.045 3.560 ;
        RECT  17.600 1.350 17.760 1.690 ;
        RECT  17.705 2.740 17.760 3.560 ;
        RECT  17.300 2.940 17.705 3.220 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.760 2.165 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.875 1.685 4.215 2.045 ;
        RECT  3.820 1.815 3.875 2.045 ;
        RECT  3.515 1.815 3.820 2.100 ;
        RECT  3.440 1.820 3.515 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 2.380 1.180 2.660 ;
        RECT  0.910 1.985 1.030 2.660 ;
        RECT  0.800 1.810 0.910 2.660 ;
        RECT  0.680 1.810 0.800 2.215 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.030 -0.400 18.480 0.400 ;
        RECT  17.510 -0.400 18.030 0.575 ;
        RECT  15.935 -0.400 17.510 0.400 ;
        RECT  15.595 -0.400 15.935 0.575 ;
        RECT  13.065 -0.400 15.595 0.400 ;
        RECT  11.565 -0.400 13.065 0.575 ;
        RECT  8.965 -0.400 11.565 0.400 ;
        RECT  8.625 -0.400 8.965 1.065 ;
        RECT  7.360 -0.400 8.625 0.400 ;
        RECT  7.020 -0.400 7.360 1.235 ;
        RECT  4.300 -0.400 7.020 0.400 ;
        RECT  2.380 -0.400 4.300 0.575 ;
        RECT  0.640 -0.400 2.380 0.400 ;
        RECT  0.300 -0.400 0.640 0.575 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.285 4.640 18.480 5.440 ;
        RECT  16.945 4.465 17.285 5.440 ;
        RECT  14.380 4.640 16.945 5.440 ;
        RECT  14.040 4.465 14.380 5.440 ;
        RECT  8.655 4.640 14.040 5.440 ;
        RECT  7.335 4.465 8.655 5.440 ;
        RECT  4.075 4.640 7.335 5.440 ;
        RECT  3.735 4.465 4.075 5.440 ;
        RECT  1.025 4.640 3.735 5.440 ;
        RECT  0.795 3.795 1.025 5.440 ;
        RECT  0.000 4.640 0.795 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.995 2.030 17.530 2.370 ;
        RECT  16.945 2.030 16.995 4.175 ;
        RECT  16.765 1.460 16.945 4.175 ;
        RECT  16.715 1.460 16.765 2.260 ;
        RECT  16.510 3.945 16.765 4.175 ;
        RECT  16.170 3.945 16.510 4.370 ;
        RECT  13.655 3.945 16.170 4.175 ;
        RECT  15.520 1.650 15.750 3.615 ;
        RECT  15.020 1.650 15.520 1.880 ;
        RECT  15.160 3.385 15.520 3.615 ;
        RECT  13.915 2.600 15.130 2.830 ;
        RECT  14.625 1.190 15.020 1.880 ;
        RECT  13.805 0.635 14.690 0.865 ;
        RECT  13.820 1.650 14.625 1.880 ;
        RECT  13.685 2.550 13.915 3.710 ;
        RECT  13.590 1.650 13.820 2.030 ;
        RECT  13.575 0.635 13.805 1.040 ;
        RECT  13.355 2.550 13.685 2.780 ;
        RECT  13.190 3.480 13.685 3.710 ;
        RECT  13.425 3.945 13.655 4.355 ;
        RECT  11.320 0.810 13.575 1.040 ;
        RECT  9.115 4.125 13.425 4.355 ;
        RECT  13.125 1.275 13.355 2.780 ;
        RECT  12.890 3.015 13.300 3.245 ;
        RECT  12.960 3.480 13.190 3.865 ;
        RECT  12.435 1.275 13.125 1.505 ;
        RECT  12.680 3.635 12.960 3.865 ;
        RECT  12.660 1.805 12.890 3.245 ;
        RECT  12.090 1.805 12.660 2.035 ;
        RECT  12.195 2.425 12.425 3.835 ;
        RECT  9.575 3.605 12.195 3.835 ;
        RECT  11.860 1.535 12.090 2.035 ;
        RECT  10.845 1.535 11.860 1.765 ;
        RECT  11.525 2.800 11.755 3.315 ;
        RECT  10.040 3.085 11.525 3.315 ;
        RECT  11.090 0.630 11.320 1.040 ;
        RECT  9.710 0.630 11.090 0.860 ;
        RECT  10.730 1.095 10.845 1.765 ;
        RECT  10.730 2.625 10.840 2.855 ;
        RECT  10.500 1.095 10.730 2.855 ;
        RECT  10.475 1.095 10.500 1.875 ;
        RECT  10.000 1.535 10.475 1.875 ;
        RECT  9.810 3.075 10.040 3.315 ;
        RECT  8.630 2.445 9.920 2.675 ;
        RECT  7.945 3.075 9.810 3.305 ;
        RECT  9.480 0.630 9.710 1.525 ;
        RECT  9.345 3.540 9.575 3.835 ;
        RECT  8.630 1.295 9.480 1.525 ;
        RECT  6.605 3.540 9.345 3.770 ;
        RECT  8.885 4.005 9.115 4.355 ;
        RECT  7.095 4.005 8.885 4.235 ;
        RECT  8.400 1.295 8.630 2.675 ;
        RECT  8.290 1.735 8.400 2.075 ;
        RECT  8.055 1.000 8.165 1.340 ;
        RECT  7.945 1.000 8.055 2.495 ;
        RECT  7.825 1.000 7.945 3.305 ;
        RECT  7.660 2.265 7.825 3.305 ;
        RECT  6.740 2.265 7.660 2.495 ;
        RECT  6.080 1.595 7.510 1.825 ;
        RECT  6.865 4.005 7.095 4.410 ;
        RECT  4.785 4.180 6.865 4.410 ;
        RECT  6.375 3.540 6.605 3.950 ;
        RECT  5.380 3.720 6.375 3.950 ;
        RECT  5.850 1.010 6.080 3.470 ;
        RECT  5.655 1.010 5.850 1.350 ;
        RECT  5.150 1.555 5.380 3.950 ;
        RECT  3.220 1.015 5.190 1.245 ;
        RECT  5.055 1.555 5.150 1.900 ;
        RECT  2.805 2.835 5.150 3.065 ;
        RECT  5.000 1.560 5.055 1.900 ;
        RECT  2.625 2.335 4.920 2.565 ;
        RECT  4.555 3.875 4.785 4.410 ;
        RECT  3.035 3.310 4.775 3.540 ;
        RECT  1.280 3.875 4.555 4.105 ;
        RECT  2.880 1.015 3.220 1.380 ;
        RECT  2.575 2.835 2.805 3.560 ;
        RECT  2.395 1.250 2.625 2.565 ;
        RECT  0.465 3.330 2.575 3.560 ;
        RECT  1.920 1.250 2.395 1.480 ;
        RECT  2.345 2.335 2.395 2.565 ;
        RECT  2.115 2.335 2.345 3.100 ;
        RECT  1.580 1.140 1.920 1.480 ;
        RECT  0.440 1.140 0.520 1.480 ;
        RECT  0.440 2.810 0.465 3.560 ;
        RECT  0.210 1.140 0.440 3.560 ;
        RECT  0.180 1.140 0.210 1.480 ;
    END
END JKFFRX1

MACRO JKFFXL
    CLASS CORE ;
    FOREIGN JKFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.780 0.810 13.010 3.755 ;
        RECT  12.680 0.810 12.780 1.285 ;
        RECT  12.400 3.525 12.780 3.755 ;
        RECT  12.405 0.810 12.680 1.040 ;
        RECT  12.175 0.730 12.405 1.040 ;
        RECT  12.060 3.525 12.400 4.190 ;
        RECT  12.030 0.730 12.175 0.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.615 1.220 13.670 1.560 ;
        RECT  13.605 2.890 13.660 3.450 ;
        RECT  13.615 1.845 13.645 2.075 ;
        RECT  13.605 1.220 13.615 2.075 ;
        RECT  13.385 1.220 13.605 3.450 ;
        RECT  13.330 1.220 13.385 1.560 ;
        RECT  13.375 1.845 13.385 3.450 ;
        RECT  13.320 2.890 13.375 3.450 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.785 3.770 2.165 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 3.490 1.120 3.910 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 1.935 2.070 2.165 ;
        RECT  1.385 1.770 1.790 2.165 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.110 -0.400 13.860 0.400 ;
        RECT  12.770 -0.400 13.110 0.575 ;
        RECT  11.610 -0.400 12.770 0.400 ;
        RECT  11.270 -0.400 11.610 1.485 ;
        RECT  8.970 -0.400 11.270 0.400 ;
        RECT  8.630 -0.400 8.970 1.400 ;
        RECT  6.600 -0.400 8.630 0.400 ;
        RECT  6.260 -0.400 6.600 0.575 ;
        RECT  3.180 -0.400 6.260 0.400 ;
        RECT  2.840 -0.400 3.180 0.575 ;
        RECT  1.680 -0.400 2.840 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.100 4.640 13.860 5.440 ;
        RECT  12.760 4.465 13.100 5.440 ;
        RECT  11.640 4.640 12.760 5.440 ;
        RECT  11.300 4.465 11.640 5.440 ;
        RECT  8.380 4.640 11.300 5.440 ;
        RECT  8.040 3.760 8.380 5.440 ;
        RECT  6.865 4.640 8.040 5.440 ;
        RECT  6.635 4.115 6.865 5.440 ;
        RECT  3.925 4.640 6.635 5.440 ;
        RECT  3.695 3.800 3.925 5.440 ;
        RECT  1.865 4.640 3.695 5.440 ;
        RECT  1.635 3.770 1.865 5.440 ;
        RECT  0.520 4.640 1.635 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.415 2.050 12.535 3.180 ;
        RECT  12.410 1.520 12.415 3.180 ;
        RECT  12.305 1.440 12.410 3.180 ;
        RECT  12.185 1.440 12.305 2.335 ;
        RECT  12.060 2.820 12.305 3.180 ;
        RECT  12.070 1.440 12.185 1.780 ;
        RECT  11.700 2.950 12.060 3.180 ;
        RECT  10.590 2.050 11.910 2.390 ;
        RECT  11.470 2.950 11.700 3.935 ;
        RECT  10.970 3.705 11.470 3.935 ;
        RECT  10.300 3.650 10.640 3.990 ;
        RECT  10.570 2.050 10.590 3.310 ;
        RECT  10.360 1.170 10.570 3.310 ;
        RECT  10.340 1.170 10.360 2.280 ;
        RECT  10.310 3.080 10.360 3.310 ;
        RECT  10.250 1.170 10.340 1.400 ;
        RECT  9.970 3.080 10.310 3.420 ;
        RECT  9.700 3.650 10.300 3.880 ;
        RECT  9.910 1.060 10.250 1.400 ;
        RECT  9.700 1.860 9.990 2.200 ;
        RECT  9.470 1.735 9.700 3.880 ;
        RECT  8.240 1.735 9.470 1.965 ;
        RECT  8.040 2.925 9.470 3.155 ;
        RECT  7.160 2.255 9.230 2.485 ;
        RECT  7.990 1.115 8.240 1.965 ;
        RECT  7.975 1.115 7.990 1.345 ;
        RECT  7.745 0.835 7.975 1.345 ;
        RECT  7.530 3.745 7.770 3.975 ;
        RECT  5.300 0.835 7.745 1.065 ;
        RECT  7.160 3.195 7.580 3.425 ;
        RECT  7.300 3.655 7.530 3.975 ;
        RECT  6.105 3.655 7.300 3.885 ;
        RECT  7.145 1.440 7.160 3.425 ;
        RECT  6.930 1.310 7.145 3.425 ;
        RECT  6.915 1.310 6.930 1.670 ;
        RECT  6.270 2.590 6.930 2.930 ;
        RECT  5.645 1.910 6.695 2.260 ;
        RECT  5.875 3.655 6.105 4.195 ;
        RECT  5.185 3.965 5.875 4.195 ;
        RECT  5.415 1.365 5.645 3.680 ;
        RECT  4.900 1.365 5.415 1.595 ;
        RECT  4.955 2.880 5.185 4.195 ;
        RECT  4.820 2.880 4.955 3.110 ;
        RECT  4.820 1.940 4.930 2.280 ;
        RECT  4.670 1.940 4.820 3.110 ;
        RECT  4.495 3.340 4.725 3.860 ;
        RECT  4.590 0.840 4.670 3.110 ;
        RECT  4.440 0.840 4.590 2.170 ;
        RECT  2.140 2.875 4.590 3.105 ;
        RECT  3.060 3.340 4.495 3.570 ;
        RECT  2.480 0.840 4.440 1.070 ;
        RECT  4.125 2.415 4.260 2.645 ;
        RECT  3.895 2.395 4.125 2.645 ;
        RECT  1.120 2.395 3.895 2.625 ;
        RECT  2.560 1.310 3.880 1.540 ;
        RECT  2.830 3.340 3.060 3.930 ;
        RECT  2.620 3.700 2.830 3.930 ;
        RECT  2.280 3.700 2.620 4.040 ;
        RECT  2.330 1.310 2.560 1.580 ;
        RECT  2.250 0.630 2.480 1.070 ;
        RECT  2.180 1.350 2.330 1.580 ;
        RECT  2.140 0.630 2.250 0.860 ;
        RECT  0.890 2.395 1.120 3.170 ;
        RECT  0.780 2.420 0.890 3.170 ;
        RECT  0.520 2.420 0.780 2.650 ;
        RECT  0.290 1.320 0.520 2.650 ;
        RECT  0.180 1.320 0.290 1.660 ;
    END
END JKFFXL

MACRO JKFFX4
    CLASS CORE ;
    FOREIGN JKFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.640 1.260 17.680 2.660 ;
        RECT  17.220 1.260 17.640 3.065 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.600 1.260 19.020 3.065 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 1.820 4.225 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.090 1.820 3.050 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 1.820 1.170 2.280 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 -0.400 19.800 0.400 ;
        RECT  19.280 -0.400 19.620 0.950 ;
        RECT  18.295 -0.400 19.280 0.400 ;
        RECT  17.955 -0.400 18.295 0.950 ;
        RECT  16.950 -0.400 17.955 0.400 ;
        RECT  16.610 -0.400 16.950 0.950 ;
        RECT  15.470 -0.400 16.610 0.400 ;
        RECT  15.130 -0.400 15.470 0.575 ;
        RECT  12.265 -0.400 15.130 0.400 ;
        RECT  11.925 -0.400 12.265 0.575 ;
        RECT  9.470 -0.400 11.925 0.400 ;
        RECT  9.130 -0.400 9.470 1.230 ;
        RECT  7.250 -0.400 9.130 0.400 ;
        RECT  6.910 -0.400 7.250 0.575 ;
        RECT  3.875 -0.400 6.910 0.400 ;
        RECT  3.535 -0.400 3.875 0.575 ;
        RECT  1.155 -0.400 3.535 0.400 ;
        RECT  0.815 -0.400 1.155 0.575 ;
        RECT  0.000 -0.400 0.815 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 4.640 19.800 5.440 ;
        RECT  19.280 3.860 19.620 5.440 ;
        RECT  18.295 4.640 19.280 5.440 ;
        RECT  17.955 3.860 18.295 5.440 ;
        RECT  16.920 4.640 17.955 5.440 ;
        RECT  16.580 4.465 16.920 5.440 ;
        RECT  15.640 4.640 16.580 5.440 ;
        RECT  15.300 4.465 15.640 5.440 ;
        RECT  13.145 4.640 15.300 5.440 ;
        RECT  12.805 4.145 13.145 5.440 ;
        RECT  10.500 4.640 12.805 5.440 ;
        RECT  9.560 4.465 10.500 5.440 ;
        RECT  7.725 4.640 9.560 5.440 ;
        RECT  7.385 4.465 7.725 5.440 ;
        RECT  4.530 4.640 7.385 5.440 ;
        RECT  4.190 4.465 4.530 5.440 ;
        RECT  2.450 4.640 4.190 5.440 ;
        RECT  2.070 4.465 2.450 5.440 ;
        RECT  1.150 4.640 2.070 5.440 ;
        RECT  0.810 4.040 1.150 5.440 ;
        RECT  0.000 4.640 0.810 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.535 2.210 19.590 2.550 ;
        RECT  19.305 2.210 19.535 3.585 ;
        RECT  19.250 2.210 19.305 2.550 ;
        RECT  16.955 3.355 19.305 3.585 ;
        RECT  16.725 1.240 16.955 3.585 ;
        RECT  16.230 1.240 16.725 1.470 ;
        RECT  16.270 2.805 16.725 3.035 ;
        RECT  16.110 2.020 16.450 2.360 ;
        RECT  16.160 2.750 16.270 3.090 ;
        RECT  16.000 0.870 16.230 1.470 ;
        RECT  15.930 2.750 16.160 3.915 ;
        RECT  15.445 2.075 16.110 2.305 ;
        RECT  15.890 0.870 16.000 1.210 ;
        RECT  15.180 3.685 15.930 3.915 ;
        RECT  15.215 1.170 15.445 3.390 ;
        RECT  13.760 1.170 15.215 1.400 ;
        RECT  14.350 3.160 15.215 3.390 ;
        RECT  14.840 3.685 15.180 4.120 ;
        RECT  12.470 3.685 14.840 3.915 ;
        RECT  14.685 2.420 14.740 2.760 ;
        RECT  14.455 1.855 14.685 2.760 ;
        RECT  13.520 1.855 14.455 2.085 ;
        RECT  14.400 2.420 14.455 2.760 ;
        RECT  14.010 3.105 14.350 3.445 ;
        RECT  13.670 2.480 14.010 2.820 ;
        RECT  11.940 3.170 14.010 3.400 ;
        RECT  13.420 1.060 13.760 1.400 ;
        RECT  12.240 2.535 13.670 2.765 ;
        RECT  13.180 1.800 13.520 2.140 ;
        RECT  12.305 1.060 13.420 1.290 ;
        RECT  10.510 1.855 13.180 2.085 ;
        RECT  12.240 3.685 12.470 4.175 ;
        RECT  12.075 1.000 12.305 1.290 ;
        RECT  11.900 2.480 12.240 2.820 ;
        RECT  7.155 3.945 12.240 4.175 ;
        RECT  10.875 1.000 12.075 1.230 ;
        RECT  11.600 3.170 11.940 3.510 ;
        RECT  11.095 2.535 11.900 2.765 ;
        RECT  10.865 2.535 11.095 3.585 ;
        RECT  10.535 0.890 10.875 1.230 ;
        RECT  8.910 3.355 10.865 3.585 ;
        RECT  10.475 1.720 10.510 2.085 ;
        RECT  10.400 1.545 10.475 2.085 ;
        RECT  10.170 1.545 10.400 3.020 ;
        RECT  8.750 1.545 10.170 1.775 ;
        RECT  9.745 2.790 10.170 3.020 ;
        RECT  9.785 2.090 9.840 2.430 ;
        RECT  9.500 2.090 9.785 2.455 ;
        RECT  9.395 2.790 9.745 3.075 ;
        RECT  8.450 2.225 9.500 2.455 ;
        RECT  8.560 3.355 8.910 3.640 ;
        RECT  8.640 0.900 8.750 1.775 ;
        RECT  8.520 0.865 8.640 1.775 ;
        RECT  6.695 3.355 8.560 3.585 ;
        RECT  8.410 0.865 8.520 1.240 ;
        RECT  8.110 2.225 8.450 3.085 ;
        RECT  6.445 0.865 8.410 1.095 ;
        RECT  8.065 2.225 8.110 2.575 ;
        RECT  7.835 1.385 8.065 2.575 ;
        RECT  7.695 1.385 7.835 1.685 ;
        RECT  7.245 2.345 7.835 2.575 ;
        RECT  7.040 1.640 7.380 1.980 ;
        RECT  6.960 2.345 7.245 2.690 ;
        RECT  6.925 3.945 7.155 4.365 ;
        RECT  6.235 1.695 7.040 1.925 ;
        RECT  6.905 2.350 6.960 2.690 ;
        RECT  5.225 4.135 6.925 4.365 ;
        RECT  6.465 3.355 6.695 3.880 ;
        RECT  6.330 3.595 6.465 3.880 ;
        RECT  6.220 0.740 6.445 1.095 ;
        RECT  5.720 3.595 6.330 3.825 ;
        RECT  6.005 1.390 6.235 3.305 ;
        RECT  6.215 0.685 6.220 1.095 ;
        RECT  5.870 0.685 6.215 0.970 ;
        RECT  5.865 1.390 6.005 1.620 ;
        RECT  5.950 2.920 6.005 3.305 ;
        RECT  5.525 1.280 5.865 1.620 ;
        RECT  5.570 2.795 5.720 3.825 ;
        RECT  5.570 1.900 5.625 2.240 ;
        RECT  5.490 1.900 5.570 3.825 ;
        RECT  5.340 1.900 5.490 3.025 ;
        RECT  5.285 1.900 5.340 2.240 ;
        RECT  2.575 2.795 5.340 3.025 ;
        RECT  4.920 3.365 5.260 3.705 ;
        RECT  4.995 3.945 5.225 4.365 ;
        RECT  3.510 3.945 4.995 4.175 ;
        RECT  4.890 2.055 4.945 2.395 ;
        RECT  3.150 3.420 4.920 3.650 ;
        RECT  4.605 2.055 4.890 2.560 ;
        RECT  2.030 2.330 4.605 2.560 ;
        RECT  4.245 1.230 4.585 1.570 ;
        RECT  3.170 1.285 4.245 1.515 ;
        RECT  3.170 3.945 3.510 4.360 ;
        RECT  2.830 1.220 3.170 1.560 ;
        RECT  1.780 3.945 3.170 4.175 ;
        RECT  2.810 3.365 3.150 3.705 ;
        RECT  2.345 2.795 2.575 3.580 ;
        RECT  2.130 1.245 2.470 1.585 ;
        RECT  0.540 3.350 2.345 3.580 ;
        RECT  1.815 1.355 2.130 1.585 ;
        RECT  1.815 2.330 2.030 3.100 ;
        RECT  1.690 1.355 1.815 3.100 ;
        RECT  1.440 3.890 1.780 4.230 ;
        RECT  1.585 1.355 1.690 2.560 ;
        RECT  0.415 2.880 0.540 3.580 ;
        RECT  0.415 1.205 0.485 1.570 ;
        RECT  0.310 1.205 0.415 3.580 ;
        RECT  0.200 1.205 0.310 3.220 ;
        RECT  0.185 1.205 0.200 3.165 ;
    END
END JKFFX4

MACRO JKFFX2
    CLASS CORE ;
    FOREIGN JKFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.855 1.755 15.085 3.195 ;
        RECT  14.830 1.755 14.855 1.985 ;
        RECT  14.735 2.635 14.855 3.195 ;
        RECT  14.600 0.640 14.830 1.985 ;
        RECT  14.700 2.635 14.735 3.080 ;
        RECT  14.490 0.640 14.600 1.450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.270 1.375 16.360 4.340 ;
        RECT  16.130 0.795 16.270 4.340 ;
        RECT  15.930 0.795 16.130 1.605 ;
        RECT  15.980 2.740 16.130 4.340 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.090 1.770 3.770 2.150 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.730 1.105 4.315 ;
        RECT  0.600 3.730 0.875 4.070 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 2.010 1.990 2.360 ;
        RECT  1.535 1.845 1.765 2.360 ;
        RECT  1.485 2.010 1.535 2.360 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.550 -0.400 16.500 0.400 ;
        RECT  15.210 -0.400 15.550 1.475 ;
        RECT  13.370 -0.400 15.210 0.400 ;
        RECT  13.030 -0.400 13.370 0.575 ;
        RECT  11.385 -0.400 13.030 0.400 ;
        RECT  11.045 -0.400 11.385 0.990 ;
        RECT  8.590 -0.400 11.045 0.400 ;
        RECT  8.250 -0.400 8.590 0.575 ;
        RECT  6.500 -0.400 8.250 0.400 ;
        RECT  6.160 -0.400 6.500 0.575 ;
        RECT  3.180 -0.400 6.160 0.400 ;
        RECT  2.840 -0.400 3.180 0.575 ;
        RECT  1.680 -0.400 2.840 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.680 4.640 16.500 5.440 ;
        RECT  15.340 4.050 15.680 5.440 ;
        RECT  13.780 4.640 15.340 5.440 ;
        RECT  13.440 4.465 13.780 5.440 ;
        RECT  11.710 4.640 13.440 5.440 ;
        RECT  11.370 3.770 11.710 5.440 ;
        RECT  8.755 4.640 11.370 5.440 ;
        RECT  8.415 3.845 8.755 5.440 ;
        RECT  6.725 4.640 8.415 5.440 ;
        RECT  6.495 4.115 6.725 5.440 ;
        RECT  3.885 4.640 6.495 5.440 ;
        RECT  3.885 3.825 3.945 4.055 ;
        RECT  3.655 3.825 3.885 5.440 ;
        RECT  3.600 3.825 3.655 4.055 ;
        RECT  1.865 4.640 3.655 5.440 ;
        RECT  1.635 4.090 1.865 5.440 ;
        RECT  0.520 4.640 1.635 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.750 1.985 15.895 2.375 ;
        RECT  15.665 1.985 15.750 3.730 ;
        RECT  15.520 2.145 15.665 3.730 ;
        RECT  14.340 3.500 15.520 3.730 ;
        RECT  14.300 3.005 14.340 3.815 ;
        RECT  14.230 1.695 14.300 3.815 ;
        RECT  14.130 1.695 14.230 3.935 ;
        RECT  14.070 1.330 14.130 3.935 ;
        RECT  13.900 1.330 14.070 1.925 ;
        RECT  14.000 3.005 14.070 3.935 ;
        RECT  12.910 3.705 14.000 3.935 ;
        RECT  13.790 1.330 13.900 1.670 ;
        RECT  13.560 2.170 13.840 2.510 ;
        RECT  13.500 1.440 13.560 2.510 ;
        RECT  13.330 1.440 13.500 2.455 ;
        RECT  12.210 1.440 13.330 1.670 ;
        RECT  13.195 2.225 13.330 2.455 ;
        RECT  12.965 2.225 13.195 3.260 ;
        RECT  12.410 3.030 12.965 3.260 ;
        RECT  12.475 2.375 12.620 2.605 ;
        RECT  12.245 1.900 12.475 2.605 ;
        RECT  12.180 3.030 12.410 3.995 ;
        RECT  10.065 1.900 12.245 2.130 ;
        RECT  11.870 1.330 12.210 1.670 ;
        RECT  12.005 3.265 12.180 3.995 ;
        RECT  11.090 3.265 12.005 3.495 ;
        RECT  10.705 2.365 11.950 2.595 ;
        RECT  10.635 1.330 11.870 1.560 ;
        RECT  10.860 3.265 11.090 4.000 ;
        RECT  10.090 3.770 10.860 4.000 ;
        RECT  10.525 2.365 10.705 2.910 ;
        RECT  10.405 1.030 10.635 1.560 ;
        RECT  10.475 2.365 10.525 3.445 ;
        RECT  10.295 2.680 10.475 3.445 ;
        RECT  10.100 1.030 10.405 1.260 ;
        RECT  9.315 3.215 10.295 3.445 ;
        RECT  9.760 0.920 10.100 1.260 ;
        RECT  9.945 1.630 10.065 2.130 ;
        RECT  9.715 1.630 9.945 2.980 ;
        RECT  9.660 1.630 9.715 1.860 ;
        RECT  8.415 2.750 9.715 2.980 ;
        RECT  9.320 1.520 9.660 1.860 ;
        RECT  7.280 2.255 9.480 2.485 ;
        RECT  7.845 1.630 9.320 1.860 ;
        RECT  9.085 3.215 9.315 3.615 ;
        RECT  8.165 3.385 9.085 3.615 ;
        RECT  8.185 2.750 8.415 3.155 ;
        RECT  8.040 2.925 8.185 3.155 ;
        RECT  7.935 3.385 8.165 4.265 ;
        RECT  7.530 4.035 7.935 4.265 ;
        RECT  7.615 0.835 7.845 1.860 ;
        RECT  5.300 0.835 7.615 1.065 ;
        RECT  7.280 3.195 7.540 3.425 ;
        RECT  7.300 3.655 7.530 4.265 ;
        RECT  6.105 3.655 7.300 3.885 ;
        RECT  7.160 2.255 7.280 3.425 ;
        RECT  7.145 1.440 7.160 3.425 ;
        RECT  6.930 1.310 7.145 3.425 ;
        RECT  6.915 1.310 6.930 1.670 ;
        RECT  6.270 2.590 6.930 2.930 ;
        RECT  5.645 1.910 6.695 2.260 ;
        RECT  5.875 3.655 6.105 4.195 ;
        RECT  5.145 3.965 5.875 4.195 ;
        RECT  5.605 1.365 5.645 2.260 ;
        RECT  5.415 1.365 5.605 3.680 ;
        RECT  4.900 1.365 5.415 1.595 ;
        RECT  5.375 2.030 5.415 3.680 ;
        RECT  4.915 2.880 5.145 4.195 ;
        RECT  4.820 1.940 4.950 2.280 ;
        RECT  4.820 2.880 4.915 3.110 ;
        RECT  4.670 1.940 4.820 3.110 ;
        RECT  4.455 3.340 4.685 3.860 ;
        RECT  4.590 0.840 4.670 3.110 ;
        RECT  4.440 0.840 4.590 2.170 ;
        RECT  2.910 2.880 4.590 3.110 ;
        RECT  3.370 3.340 4.455 3.570 ;
        RECT  2.440 0.840 4.440 1.070 ;
        RECT  2.450 2.420 4.280 2.650 ;
        RECT  2.560 1.310 3.880 1.540 ;
        RECT  3.140 3.340 3.370 4.345 ;
        RECT  2.280 4.115 3.140 4.345 ;
        RECT  2.680 2.880 2.910 3.315 ;
        RECT  2.140 3.085 2.680 3.315 ;
        RECT  2.330 1.310 2.560 1.745 ;
        RECT  2.220 2.420 2.450 2.855 ;
        RECT  2.100 0.630 2.440 1.070 ;
        RECT  2.140 1.515 2.330 1.745 ;
        RECT  1.065 2.625 2.220 2.855 ;
        RECT  0.835 2.420 1.065 3.375 ;
        RECT  0.520 2.420 0.835 2.650 ;
        RECT  0.290 1.350 0.520 2.650 ;
        RECT  0.180 1.350 0.290 1.690 ;
    END
END JKFFX2

MACRO JKFFX1
    CLASS CORE ;
    FOREIGN JKFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.765 0.810 12.995 3.755 ;
        RECT  12.425 0.810 12.765 1.040 ;
        RECT  12.400 3.525 12.765 3.755 ;
        RECT  12.195 0.745 12.425 1.040 ;
        RECT  12.095 3.525 12.400 4.030 ;
        RECT  12.050 0.745 12.195 0.975 ;
        RECT  12.060 3.690 12.095 4.030 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 1.820 13.720 3.220 ;
        RECT  13.650 1.820 13.660 3.570 ;
        RECT  13.340 1.300 13.650 3.570 ;
        RECT  13.310 1.300 13.340 1.640 ;
        RECT  13.320 2.760 13.340 3.570 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.770 3.770 2.150 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 3.490 1.120 3.910 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 1.935 2.070 2.165 ;
        RECT  1.385 1.770 1.790 2.165 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.090 -0.400 13.860 0.400 ;
        RECT  12.750 -0.400 13.090 0.575 ;
        RECT  11.630 -0.400 12.750 0.400 ;
        RECT  11.290 -0.400 11.630 1.420 ;
        RECT  8.990 -0.400 11.290 0.400 ;
        RECT  8.650 -0.400 8.990 1.280 ;
        RECT  6.500 -0.400 8.650 0.400 ;
        RECT  6.160 -0.400 6.500 0.575 ;
        RECT  3.180 -0.400 6.160 0.400 ;
        RECT  2.840 -0.400 3.180 0.575 ;
        RECT  1.680 -0.400 2.840 0.400 ;
        RECT  1.340 -0.400 1.680 0.575 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.940 4.640 13.860 5.440 ;
        RECT  12.600 4.465 12.940 5.440 ;
        RECT  11.640 4.640 12.600 5.440 ;
        RECT  11.300 4.465 11.640 5.440 ;
        RECT  8.380 4.640 11.300 5.440 ;
        RECT  8.040 3.760 8.380 5.440 ;
        RECT  6.865 4.640 8.040 5.440 ;
        RECT  6.635 4.115 6.865 5.440 ;
        RECT  3.925 4.640 6.635 5.440 ;
        RECT  3.695 3.800 3.925 5.440 ;
        RECT  1.865 4.640 3.695 5.440 ;
        RECT  1.635 3.770 1.865 5.440 ;
        RECT  0.520 4.640 1.635 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.390 1.520 12.535 3.180 ;
        RECT  12.305 1.460 12.390 3.180 ;
        RECT  12.050 1.460 12.305 1.800 ;
        RECT  12.060 2.840 12.305 3.180 ;
        RECT  11.700 2.950 12.060 3.180 ;
        RECT  10.590 2.050 11.910 2.390 ;
        RECT  11.470 2.950 11.700 3.935 ;
        RECT  10.970 3.705 11.470 3.935 ;
        RECT  10.300 3.650 10.640 3.990 ;
        RECT  10.360 1.170 10.590 3.170 ;
        RECT  10.270 1.170 10.360 1.400 ;
        RECT  10.270 2.940 10.360 3.170 ;
        RECT  9.700 3.650 10.300 3.880 ;
        RECT  9.930 1.060 10.270 1.400 ;
        RECT  9.930 2.940 10.270 3.280 ;
        RECT  9.700 1.860 10.010 2.200 ;
        RECT  9.470 1.735 9.700 3.880 ;
        RECT  8.240 1.735 9.470 1.965 ;
        RECT  8.040 2.925 9.470 3.155 ;
        RECT  7.160 2.255 9.240 2.485 ;
        RECT  8.010 0.985 8.240 1.965 ;
        RECT  7.975 0.985 8.010 1.215 ;
        RECT  7.745 0.835 7.975 1.215 ;
        RECT  7.530 3.745 7.770 3.975 ;
        RECT  5.300 0.835 7.745 1.065 ;
        RECT  7.160 3.195 7.580 3.425 ;
        RECT  7.300 3.655 7.530 3.975 ;
        RECT  6.105 3.655 7.300 3.885 ;
        RECT  7.145 1.440 7.160 3.425 ;
        RECT  6.930 1.310 7.145 3.425 ;
        RECT  6.915 1.310 6.930 1.670 ;
        RECT  6.270 2.590 6.930 2.930 ;
        RECT  5.645 1.910 6.695 2.260 ;
        RECT  5.875 3.655 6.105 4.195 ;
        RECT  5.185 3.965 5.875 4.195 ;
        RECT  5.415 1.365 5.645 3.680 ;
        RECT  4.900 1.365 5.415 1.595 ;
        RECT  4.955 2.880 5.185 4.195 ;
        RECT  4.820 2.880 4.955 3.110 ;
        RECT  4.820 1.940 4.930 2.280 ;
        RECT  4.670 1.940 4.820 3.110 ;
        RECT  4.495 3.340 4.725 3.860 ;
        RECT  4.590 0.840 4.670 3.110 ;
        RECT  4.440 0.840 4.590 2.170 ;
        RECT  2.140 2.880 4.590 3.110 ;
        RECT  3.060 3.340 4.495 3.570 ;
        RECT  2.440 0.840 4.440 1.070 ;
        RECT  1.120 2.420 4.260 2.650 ;
        RECT  2.560 1.310 3.880 1.540 ;
        RECT  2.830 3.340 3.060 3.930 ;
        RECT  2.620 3.700 2.830 3.930 ;
        RECT  2.280 3.700 2.620 4.040 ;
        RECT  2.330 1.310 2.560 1.635 ;
        RECT  2.155 0.630 2.440 1.070 ;
        RECT  2.140 1.405 2.330 1.635 ;
        RECT  2.100 0.630 2.155 0.970 ;
        RECT  0.780 2.420 1.120 3.170 ;
        RECT  0.520 2.420 0.780 2.650 ;
        RECT  0.290 1.350 0.520 2.650 ;
        RECT  0.180 1.350 0.290 1.690 ;
    END
END JKFFX1

MACRO INVXL
    CLASS CORE ;
    FOREIGN INVXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 2.380 1.180 3.225 ;
        RECT  1.030 1.350 1.120 1.845 ;
        RECT  0.800 1.350 1.030 3.225 ;
        RECT  0.780 1.350 0.800 1.845 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.520 2.510 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.990 -0.400 1.320 0.400 ;
        RECT  0.180 -0.400 0.990 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.850 4.640 1.320 5.440 ;
        RECT  0.850 3.820 1.085 4.160 ;
        RECT  0.510 3.820 0.850 5.440 ;
        RECT  0.275 3.820 0.510 4.160 ;
        RECT  0.000 4.640 0.510 5.440 ;
        END
    END VDD
END INVXL

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 1.760 3.745 3.220 ;
        RECT  3.085 1.515 3.160 3.220 ;
        RECT  2.920 1.515 3.085 3.275 ;
        RECT  2.195 1.290 2.920 3.410 ;
        RECT  2.120 1.290 2.195 1.820 ;
        RECT  0.780 2.930 2.195 3.410 ;
        RECT  0.780 1.290 2.120 1.770 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.045 1.355 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 -0.400 3.960 0.400 ;
        RECT  2.945 -0.400 3.755 0.575 ;
        RECT  1.920 -0.400 2.945 0.400 ;
        RECT  1.580 -0.400 1.920 0.960 ;
        RECT  0.560 -0.400 1.580 0.400 ;
        RECT  0.220 -0.400 0.560 0.575 ;
        RECT  0.000 -0.400 0.220 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 4.640 3.960 5.440 ;
        RECT  3.320 4.465 3.780 5.440 ;
        RECT  2.980 3.790 3.320 5.440 ;
        RECT  1.915 4.640 2.980 5.440 ;
        RECT  1.575 3.790 1.915 5.440 ;
        RECT  0.520 4.640 1.575 5.440 ;
        RECT  0.180 3.790 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END INVX8

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 0.815 1.285 4.240 ;
        RECT  0.800 1.820 0.945 3.220 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.875 0.520 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 -0.400 2.640 0.400 ;
        RECT  1.705 -0.400 2.045 1.625 ;
        RECT  0.520 -0.400 1.705 0.400 ;
        RECT  0.180 -0.400 0.520 1.625 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 4.640 2.640 5.440 ;
        RECT  1.705 2.960 2.045 5.440 ;
        RECT  0.520 4.640 1.705 5.440 ;
        RECT  0.180 2.960 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END INVX4

MACRO INVX3
    CLASS CORE ;
    FOREIGN INVX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.240 1.845 3.835 ;
        RECT  0.525 1.240 1.505 1.580 ;
        RECT  1.460 2.940 1.505 3.780 ;
        RECT  0.525 3.245 1.460 3.585 ;
        RECT  0.185 0.905 0.525 1.715 ;
        RECT  0.185 3.025 0.525 3.835 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.070 1.005 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 -0.400 2.640 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 4.640 2.640 5.440 ;
        RECT  0.945 4.465 1.285 5.440 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
END INVX3

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.610 0.770 1.840 3.005 ;
        RECT  1.460 0.770 1.610 1.580 ;
        RECT  1.535 2.635 1.610 3.005 ;
        RECT  1.080 2.775 1.535 3.005 ;
        RECT  0.740 2.775 1.080 3.585 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.495 1.820 1.305 2.410 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 -0.400 1.980 0.400 ;
        RECT  0.540 -0.400 0.880 1.580 ;
        RECT  0.000 -0.400 0.540 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 4.640 1.980 5.440 ;
        RECT  1.635 4.465 1.640 5.440 ;
        RECT  1.305 4.405 1.635 5.440 ;
        RECT  1.300 4.465 1.305 5.440 ;
        RECT  0.000 4.640 1.300 5.440 ;
        END
    END VDD
END INVX2

MACRO INVX20
    CLASS CORE ;
    FOREIGN INVX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.775 1.195 12.325 3.840 ;
        RECT  10.385 1.195 10.775 1.880 ;
        RECT  10.235 2.990 10.775 3.670 ;
        RECT  7.215 1.200 10.385 1.880 ;
        RECT  9.685 2.925 10.235 3.735 ;
        RECT  8.815 2.990 9.685 3.670 ;
        RECT  8.365 2.925 8.815 3.735 ;
        RECT  7.475 2.990 8.365 3.670 ;
        RECT  7.045 2.925 7.475 3.735 ;
        RECT  6.875 1.195 7.215 1.880 ;
        RECT  6.155 2.990 7.045 3.670 ;
        RECT  5.625 1.195 6.875 1.875 ;
        RECT  5.625 2.925 6.155 3.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.100 1.255 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.335 -0.400 12.540 0.400 ;
        RECT  11.995 -0.400 12.335 0.575 ;
        RECT  10.950 -0.400 11.995 0.400 ;
        RECT  10.610 -0.400 10.950 0.575 ;
        RECT  9.530 -0.400 10.610 0.400 ;
        RECT  9.190 -0.400 9.530 0.575 ;
        RECT  8.100 -0.400 9.190 0.400 ;
        RECT  7.760 -0.400 8.100 0.575 ;
        RECT  6.680 -0.400 7.760 0.400 ;
        RECT  6.340 -0.400 6.680 0.575 ;
        RECT  5.285 -0.400 6.340 0.400 ;
        RECT  4.945 -0.400 5.285 0.575 ;
        RECT  3.840 -0.400 4.945 0.400 ;
        RECT  3.500 -0.400 3.840 1.020 ;
        RECT  2.415 -0.400 3.500 0.400 ;
        RECT  2.075 -0.400 2.415 1.020 ;
        RECT  1.005 -0.400 2.075 0.400 ;
        RECT  0.665 -0.400 1.005 1.685 ;
        RECT  0.000 -0.400 0.665 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.335 4.640 12.540 5.440 ;
        RECT  11.995 4.465 12.335 5.440 ;
        RECT  10.950 4.640 11.995 5.440 ;
        RECT  10.610 4.465 10.950 5.440 ;
        RECT  9.530 4.640 10.610 5.440 ;
        RECT  9.190 4.465 9.530 5.440 ;
        RECT  8.095 4.640 9.190 5.440 ;
        RECT  7.755 4.465 8.095 5.440 ;
        RECT  6.675 4.640 7.755 5.440 ;
        RECT  6.335 4.465 6.675 5.440 ;
        RECT  5.260 4.640 6.335 5.440 ;
        RECT  4.920 4.465 5.260 5.440 ;
        RECT  3.835 4.640 4.920 5.440 ;
        RECT  3.495 4.060 3.835 5.440 ;
        RECT  2.365 4.640 3.495 5.440 ;
        RECT  2.025 4.090 2.365 5.440 ;
        RECT  1.005 4.640 2.025 5.440 ;
        RECT  0.665 3.050 1.005 5.440 ;
        RECT  0.000 4.640 0.665 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.415 2.190 10.455 2.530 ;
        RECT  4.820 2.210 5.415 2.510 ;
        RECT  4.520 1.420 4.820 3.735 ;
        RECT  2.790 1.420 4.520 1.760 ;
        RECT  2.785 2.925 4.520 3.735 ;
        RECT  2.480 2.100 4.230 2.440 ;
        RECT  1.775 2.155 2.480 2.385 ;
        RECT  1.545 1.420 1.775 3.315 ;
        RECT  1.435 1.420 1.545 1.760 ;
        RECT  1.435 2.975 1.545 3.315 ;
    END
END INVX20

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.065 2.370 1.180 3.560 ;
        RECT  0.835 1.350 1.065 3.560 ;
        RECT  0.800 2.370 0.835 3.560 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.570 2.385 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.400 1.320 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 1.320 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END INVX1

MACRO INVX16
    CLASS CORE ;
    FOREIGN INVX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 1.200 11.005 3.840 ;
        RECT  7.215 1.200 9.455 1.880 ;
        RECT  8.815 2.990 9.455 3.670 ;
        RECT  8.365 2.925 8.815 3.735 ;
        RECT  7.475 2.990 8.365 3.670 ;
        RECT  7.045 2.925 7.475 3.735 ;
        RECT  6.875 1.195 7.215 1.880 ;
        RECT  6.155 2.990 7.045 3.670 ;
        RECT  5.625 1.195 6.875 1.875 ;
        RECT  5.625 2.925 6.155 3.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.100 1.255 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.950 -0.400 11.220 0.400 ;
        RECT  10.610 -0.400 10.950 0.575 ;
        RECT  9.530 -0.400 10.610 0.400 ;
        RECT  9.190 -0.400 9.530 0.575 ;
        RECT  8.100 -0.400 9.190 0.400 ;
        RECT  7.760 -0.400 8.100 0.575 ;
        RECT  6.675 -0.400 7.760 0.400 ;
        RECT  6.335 -0.400 6.675 0.575 ;
        RECT  5.285 -0.400 6.335 0.400 ;
        RECT  4.945 -0.400 5.285 0.575 ;
        RECT  3.840 -0.400 4.945 0.400 ;
        RECT  3.500 -0.400 3.840 1.020 ;
        RECT  2.415 -0.400 3.500 0.400 ;
        RECT  2.075 -0.400 2.415 1.020 ;
        RECT  0.965 -0.400 2.075 0.400 ;
        RECT  0.625 -0.400 0.965 1.780 ;
        RECT  0.000 -0.400 0.625 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.950 4.640 11.220 5.440 ;
        RECT  10.610 4.465 10.950 5.440 ;
        RECT  9.530 4.640 10.610 5.440 ;
        RECT  9.190 4.465 9.530 5.440 ;
        RECT  8.095 4.640 9.190 5.440 ;
        RECT  7.755 4.465 8.095 5.440 ;
        RECT  6.675 4.640 7.755 5.440 ;
        RECT  6.335 4.465 6.675 5.440 ;
        RECT  5.270 4.640 6.335 5.440 ;
        RECT  4.930 4.465 5.270 5.440 ;
        RECT  3.835 4.640 4.930 5.440 ;
        RECT  3.495 4.060 3.835 5.440 ;
        RECT  2.365 4.640 3.495 5.440 ;
        RECT  2.025 4.090 2.365 5.440 ;
        RECT  0.965 4.640 2.025 5.440 ;
        RECT  0.625 3.050 0.965 5.440 ;
        RECT  0.000 4.640 0.625 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.520 2.190 9.150 2.530 ;
        RECT  4.820 2.210 5.520 2.510 ;
        RECT  4.520 1.420 4.820 3.225 ;
        RECT  2.790 1.420 4.520 1.760 ;
        RECT  4.485 2.925 4.520 3.225 ;
        RECT  4.145 2.925 4.485 3.735 ;
        RECT  2.480 2.100 4.230 2.440 ;
        RECT  3.125 2.925 4.145 3.265 ;
        RECT  2.785 2.925 3.125 3.735 ;
        RECT  1.775 2.155 2.480 2.385 ;
        RECT  1.545 1.420 1.775 3.315 ;
        RECT  1.435 1.420 1.545 1.760 ;
        RECT  1.435 2.975 1.545 3.315 ;
    END
END INVX16

MACRO INVX12
    CLASS CORE ;
    FOREIGN INVX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.200 8.365 3.840 ;
        RECT  4.310 1.200 6.815 1.880 ;
        RECT  6.740 2.630 6.815 3.840 ;
        RECT  4.305 2.840 6.740 3.840 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.130 0.860 2.470 ;
        RECT  0.445 2.240 0.520 2.470 ;
        RECT  0.215 2.240 0.445 2.635 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.390 -0.400 8.580 0.400 ;
        RECT  8.050 -0.400 8.390 0.900 ;
        RECT  6.970 -0.400 8.050 0.400 ;
        RECT  6.630 -0.400 6.970 0.900 ;
        RECT  5.535 -0.400 6.630 0.400 ;
        RECT  5.195 -0.400 5.535 0.900 ;
        RECT  2.780 -0.400 5.195 0.400 ;
        RECT  2.440 -0.400 2.780 0.575 ;
        RECT  1.395 -0.400 2.440 0.400 ;
        RECT  1.055 -0.400 1.395 1.060 ;
        RECT  0.000 -0.400 1.055 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.400 4.640 8.580 5.440 ;
        RECT  8.060 4.090 8.400 5.440 ;
        RECT  6.970 4.640 8.060 5.440 ;
        RECT  6.630 4.090 6.970 5.440 ;
        RECT  5.535 4.640 6.630 5.440 ;
        RECT  5.195 4.090 5.535 5.440 ;
        RECT  4.140 4.640 5.195 5.440 ;
        RECT  3.795 4.410 4.140 5.440 ;
        RECT  1.340 4.640 3.795 5.440 ;
        RECT  1.000 4.465 1.340 5.440 ;
        RECT  0.000 4.640 1.000 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.490 2.190 6.510 2.530 ;
        RECT  3.190 1.420 3.490 3.220 ;
        RECT  1.755 1.420 3.190 1.760 ;
        RECT  2.095 2.880 3.190 3.220 ;
        RECT  1.415 2.100 2.660 2.440 ;
        RECT  1.755 2.880 2.095 3.730 ;
        RECT  1.185 1.440 1.415 3.235 ;
        RECT  0.540 1.440 1.185 1.670 ;
        RECT  0.520 3.005 1.185 3.235 ;
        RECT  0.200 1.440 0.540 1.780 ;
        RECT  0.180 2.895 0.520 3.235 ;
    END
END INVX12

MACRO HOLDX1
    CLASS CORE ;
    FOREIGN HOLDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION INOUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 3.180 2.165 3.520 ;
        RECT  1.880 1.515 2.110 3.520 ;
        RECT  0.980 1.515 1.880 1.745 ;
        RECT  1.825 2.720 1.880 3.520 ;
        RECT  1.535 2.720 1.825 3.195 ;
        RECT  0.870 2.720 1.535 2.950 ;
        RECT  0.640 2.550 0.870 2.950 ;
        END
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 -0.400 2.640 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 4.640 2.640 5.440 ;
        RECT  1.020 4.465 1.360 5.440 ;
        RECT  0.000 4.640 1.020 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.410 2.055 1.600 2.285 ;
        RECT  0.410 0.880 0.520 1.220 ;
        RECT  0.410 3.180 0.520 3.520 ;
        RECT  0.180 0.880 0.410 3.520 ;
    END
END HOLDX1

MACRO EDFFTRXL
    CLASS CORE ;
    FOREIGN EDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 4.015 2.120 4.340 ;
        RECT  1.460 4.015 1.820 4.410 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.795 3.640 15.905 3.980 ;
        RECT  15.625 3.135 15.795 3.980 ;
        RECT  15.565 2.075 15.625 3.980 ;
        RECT  15.540 2.075 15.565 3.365 ;
        RECT  15.395 1.350 15.540 3.365 ;
        RECT  15.310 1.350 15.395 2.385 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.845 1.025 15.075 3.520 ;
        RECT  14.650 1.025 14.845 1.255 ;
        RECT  14.660 3.195 14.845 3.520 ;
        RECT  14.465 3.290 14.660 3.520 ;
        RECT  14.475 0.740 14.650 1.255 ;
        RECT  14.420 0.685 14.475 1.255 ;
        RECT  14.235 3.290 14.465 4.315 ;
        RECT  14.135 0.685 14.420 1.025 ;
        RECT  14.125 3.575 14.235 4.315 ;
        RECT  14.075 4.085 14.125 4.315 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.655 5.025 1.885 ;
        RECT  4.235 1.655 4.465 2.045 ;
        RECT  3.085 1.815 4.235 2.045 ;
        RECT  2.855 1.815 3.085 2.240 ;
        RECT  1.850 2.010 2.855 2.240 ;
        RECT  1.620 1.860 1.850 2.240 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.355 1.845 5.800 2.335 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 2.965 1.105 3.195 ;
        RECT  0.855 2.370 0.925 3.195 ;
        RECT  0.695 2.030 0.855 3.195 ;
        RECT  0.625 2.030 0.695 2.600 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.595 -0.400 16.500 0.400 ;
        RECT  15.255 -0.400 15.595 0.575 ;
        RECT  13.755 -0.400 15.255 0.400 ;
        RECT  13.415 -0.400 13.755 1.025 ;
        RECT  11.020 -0.400 13.415 0.400 ;
        RECT  10.790 -0.400 11.020 1.415 ;
        RECT  8.200 -0.400 10.790 0.400 ;
        RECT  7.860 -0.400 8.200 0.885 ;
        RECT  1.800 -0.400 7.860 0.400 ;
        RECT  1.460 -0.400 1.800 0.575 ;
        RECT  0.000 -0.400 1.460 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.185 4.640 16.500 5.440 ;
        RECT  14.845 3.755 15.185 5.440 ;
        RECT  12.910 4.640 14.845 5.440 ;
        RECT  12.680 3.310 12.910 5.440 ;
        RECT  10.270 4.640 12.680 5.440 ;
        RECT  9.930 4.465 10.270 5.440 ;
        RECT  7.740 4.640 9.930 5.440 ;
        RECT  7.400 4.465 7.740 5.440 ;
        RECT  4.170 4.640 7.400 5.440 ;
        RECT  3.830 4.465 4.170 5.440 ;
        RECT  1.185 4.640 3.830 5.440 ;
        RECT  0.845 4.465 1.185 5.440 ;
        RECT  0.000 4.640 0.845 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.460 2.200 14.615 2.560 ;
        RECT  14.460 1.495 14.515 1.835 ;
        RECT  14.390 1.495 14.460 2.560 ;
        RECT  14.175 1.495 14.390 3.060 ;
        RECT  14.160 1.550 14.175 3.060 ;
        RECT  13.605 2.830 14.160 3.060 ;
        RECT  13.590 2.010 13.930 2.350 ;
        RECT  13.605 3.320 13.690 3.660 ;
        RECT  13.375 2.830 13.605 3.660 ;
        RECT  13.415 2.010 13.590 2.240 ;
        RECT  13.185 1.765 13.415 2.240 ;
        RECT  12.405 2.830 13.375 3.060 ;
        RECT  13.350 3.320 13.375 3.660 ;
        RECT  12.410 1.765 13.185 1.995 ;
        RECT  11.785 0.705 12.765 0.935 ;
        RECT  12.255 1.285 12.410 1.995 ;
        RECT  12.175 2.830 12.405 4.235 ;
        RECT  12.025 1.285 12.255 2.510 ;
        RECT  3.275 4.005 12.175 4.235 ;
        RECT  11.735 2.280 12.025 2.510 ;
        RECT  11.555 0.705 11.785 2.040 ;
        RECT  11.505 2.280 11.735 3.755 ;
        RECT  10.560 1.810 11.555 2.040 ;
        RECT  11.260 3.525 11.505 3.755 ;
        RECT  10.890 2.635 11.250 3.005 ;
        RECT  10.560 2.635 10.890 2.865 ;
        RECT  10.330 0.675 10.560 2.865 ;
        RECT  8.675 0.675 10.330 0.905 ;
        RECT  10.105 1.610 10.330 1.975 ;
        RECT  10.075 2.635 10.330 2.865 ;
        RECT  9.615 1.135 10.100 1.365 ;
        RECT  9.845 2.635 10.075 3.115 ;
        RECT  9.385 1.135 9.615 3.650 ;
        RECT  9.285 1.135 9.385 1.560 ;
        RECT  9.225 3.310 9.385 3.650 ;
        RECT  8.995 2.610 9.150 2.975 ;
        RECT  8.740 1.580 9.005 1.810 ;
        RECT  8.765 2.195 8.995 3.635 ;
        RECT  8.740 2.195 8.765 2.425 ;
        RECT  7.965 3.405 8.765 3.635 ;
        RECT  8.510 1.580 8.740 2.425 ;
        RECT  8.445 0.675 8.675 1.345 ;
        RECT  7.210 2.835 8.535 3.065 ;
        RECT  7.925 2.195 8.510 2.425 ;
        RECT  7.465 1.115 8.445 1.345 ;
        RECT  7.695 2.060 7.925 2.425 ;
        RECT  7.235 0.685 7.465 1.345 ;
        RECT  6.510 0.685 7.235 0.915 ;
        RECT  6.980 2.065 7.210 3.635 ;
        RECT  6.970 2.065 6.980 2.295 ;
        RECT  5.985 3.405 6.980 3.635 ;
        RECT  6.740 1.145 6.970 2.295 ;
        RECT  6.260 2.750 6.740 3.095 ;
        RECT  6.280 0.685 6.510 1.630 ;
        RECT  6.260 1.400 6.280 1.630 ;
        RECT  6.030 1.400 6.260 3.095 ;
        RECT  5.820 0.665 6.050 1.105 ;
        RECT  5.115 2.765 6.030 2.995 ;
        RECT  3.045 0.665 5.820 0.895 ;
        RECT  2.710 3.445 5.440 3.675 ;
        RECT  4.885 2.765 5.115 3.215 ;
        RECT  2.245 2.985 4.885 3.215 ;
        RECT  2.805 1.125 4.745 1.355 ;
        RECT  1.785 2.520 4.320 2.750 ;
        RECT  3.045 4.005 3.275 4.390 ;
        RECT  2.880 4.160 3.045 4.390 ;
        RECT  2.575 0.665 2.805 1.355 ;
        RECT  2.480 3.445 2.710 3.860 ;
        RECT  2.340 0.665 2.575 0.895 ;
        RECT  2.015 2.985 2.245 3.690 ;
        RECT  0.465 3.460 2.015 3.690 ;
        RECT  1.390 1.385 1.920 1.615 ;
        RECT  1.555 2.480 1.785 3.130 ;
        RECT  1.390 2.480 1.555 2.710 ;
        RECT  1.160 1.385 1.390 2.710 ;
        RECT  0.395 1.200 0.520 1.540 ;
        RECT  0.395 2.855 0.465 3.690 ;
        RECT  0.235 1.200 0.395 3.690 ;
        RECT  0.180 1.200 0.235 3.170 ;
        RECT  0.165 1.255 0.180 3.170 ;
    END
END EDFFTRXL

MACRO EDFFTRX4
    CLASS CORE ;
    FOREIGN EDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFTRXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.420 3.780 1.840 4.340 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.300 1.260 20.320 2.660 ;
        RECT  19.940 1.260 20.300 3.140 ;
        RECT  19.855 1.300 19.940 1.640 ;
        RECT  19.925 2.630 19.940 3.140 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.985 1.260 19.000 2.660 ;
        RECT  18.640 1.260 18.985 3.140 ;
        RECT  18.620 1.260 18.640 2.660 ;
        RECT  18.575 1.300 18.620 1.640 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.260 1.670 5.625 2.085 ;
        RECT  5.065 1.820 5.260 2.085 ;
        RECT  3.515 1.855 5.065 2.085 ;
        RECT  2.855 1.845 3.515 2.085 ;
        RECT  1.970 1.855 2.855 2.085 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.155 4.070 6.385 4.315 ;
        RECT  5.270 4.070 6.155 4.300 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.015 1.845 1.105 2.340 ;
        RECT  0.655 1.845 1.015 2.345 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.875 -0.400 21.120 0.400 ;
        RECT  20.535 -0.400 20.875 0.575 ;
        RECT  19.555 -0.400 20.535 0.400 ;
        RECT  19.215 -0.400 19.555 1.010 ;
        RECT  18.275 -0.400 19.215 0.400 ;
        RECT  17.935 -0.400 18.275 1.010 ;
        RECT  16.925 -0.400 17.935 0.400 ;
        RECT  16.585 -0.400 16.925 0.575 ;
        RECT  14.335 -0.400 16.585 0.400 ;
        RECT  14.105 -0.400 14.335 0.950 ;
        RECT  11.825 -0.400 14.105 0.400 ;
        RECT  11.485 -0.400 11.825 0.950 ;
        RECT  10.300 -0.400 11.485 0.400 ;
        RECT  9.960 -0.400 10.300 1.225 ;
        RECT  8.860 -0.400 9.960 0.400 ;
        RECT  8.520 -0.400 8.860 1.215 ;
        RECT  2.460 -0.400 8.520 0.400 ;
        RECT  2.120 -0.400 2.460 0.575 ;
        RECT  1.200 -0.400 2.120 0.415 ;
        RECT  0.860 -0.400 1.200 0.575 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.910 4.640 21.120 5.440 ;
        RECT  20.570 4.010 20.910 5.440 ;
        RECT  19.625 4.640 20.570 5.440 ;
        RECT  19.285 4.010 19.625 5.440 ;
        RECT  18.305 4.640 19.285 5.440 ;
        RECT  17.965 4.010 18.305 5.440 ;
        RECT  16.960 4.640 17.965 5.440 ;
        RECT  16.620 4.465 16.960 5.440 ;
        RECT  14.070 4.640 16.620 5.440 ;
        RECT  13.730 4.465 14.070 5.440 ;
        RECT  11.430 4.640 13.730 5.440 ;
        RECT  11.090 4.465 11.430 5.440 ;
        RECT  8.080 4.640 11.090 5.440 ;
        RECT  7.740 4.465 8.080 5.440 ;
        RECT  4.660 4.640 7.740 5.440 ;
        RECT  4.320 3.755 4.660 5.440 ;
        RECT  2.490 4.640 4.320 5.440 ;
        RECT  2.150 3.795 2.490 5.440 ;
        RECT  1.105 4.640 2.150 5.440 ;
        RECT  0.875 3.970 1.105 5.440 ;
        RECT  0.000 4.640 0.875 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.625 2.165 20.855 3.715 ;
        RECT  18.290 3.485 20.625 3.715 ;
        RECT  18.060 1.410 18.290 3.715 ;
        RECT  17.635 1.410 18.060 1.640 ;
        RECT  17.550 2.740 18.060 3.080 ;
        RECT  17.035 1.975 17.795 2.370 ;
        RECT  17.295 1.300 17.635 1.640 ;
        RECT  17.320 2.740 17.550 4.175 ;
        RECT  16.310 3.945 17.320 4.175 ;
        RECT  16.805 1.075 17.035 3.655 ;
        RECT  15.390 1.075 16.805 1.305 ;
        RECT  12.410 3.425 16.805 3.655 ;
        RECT  16.140 1.755 16.325 3.135 ;
        RECT  16.080 3.945 16.310 4.325 ;
        RECT  16.095 1.700 16.140 3.135 ;
        RECT  15.800 1.700 16.095 2.040 ;
        RECT  15.055 2.905 16.095 3.135 ;
        RECT  15.960 4.005 16.080 4.325 ;
        RECT  7.420 4.005 15.960 4.235 ;
        RECT  15.090 1.705 15.430 2.045 ;
        RECT  15.160 1.075 15.390 1.410 ;
        RECT  13.840 1.180 15.160 1.410 ;
        RECT  13.365 1.760 15.090 1.990 ;
        RECT  14.700 2.475 15.055 3.135 ;
        RECT  12.445 2.905 14.700 3.135 ;
        RECT  12.905 2.440 14.205 2.670 ;
        RECT  13.610 0.960 13.840 1.410 ;
        RECT  13.055 0.960 13.610 1.190 ;
        RECT  13.135 1.535 13.365 1.990 ;
        RECT  12.595 1.535 13.135 1.765 ;
        RECT  12.825 0.770 13.055 1.190 ;
        RECT  12.675 1.995 12.905 2.670 ;
        RECT  11.775 1.995 12.675 2.225 ;
        RECT  12.365 1.180 12.595 1.765 ;
        RECT  12.080 2.475 12.445 3.135 ;
        RECT  11.105 1.180 12.365 1.410 ;
        RECT  11.025 2.905 12.080 3.135 ;
        RECT  11.510 1.895 11.775 2.225 ;
        RECT  11.280 1.895 11.510 2.315 ;
        RECT  10.565 2.085 11.280 2.315 ;
        RECT  11.050 0.810 11.105 1.410 ;
        RECT  10.820 0.810 11.050 1.795 ;
        RECT  10.795 2.630 11.025 3.775 ;
        RECT  10.765 0.810 10.820 1.150 ;
        RECT  10.105 1.565 10.820 1.795 ;
        RECT  8.765 3.545 10.795 3.775 ;
        RECT  10.335 2.085 10.565 3.135 ;
        RECT  9.350 2.905 10.335 3.135 ;
        RECT  9.875 1.565 10.105 2.675 ;
        RECT  9.695 2.445 9.875 2.675 ;
        RECT  9.415 0.995 9.645 1.745 ;
        RECT  9.240 0.995 9.415 1.225 ;
        RECT  9.280 1.515 9.415 1.745 ;
        RECT  9.280 2.905 9.350 3.315 ;
        RECT  9.050 1.515 9.280 3.315 ;
        RECT  8.525 1.515 9.050 1.765 ;
        RECT  8.995 3.085 9.050 3.315 ;
        RECT  8.535 2.165 8.765 3.775 ;
        RECT  8.000 2.165 8.535 2.395 ;
        RECT  8.295 1.515 8.525 1.880 ;
        RECT  7.540 2.625 8.305 2.990 ;
        RECT  7.770 0.630 8.000 2.395 ;
        RECT  6.985 0.630 7.770 0.860 ;
        RECT  7.445 1.325 7.540 3.655 ;
        RECT  7.310 1.090 7.445 3.655 ;
        RECT  7.190 4.005 7.420 4.375 ;
        RECT  7.215 1.090 7.310 1.555 ;
        RECT  6.365 3.425 7.310 3.655 ;
        RECT  6.920 4.145 7.190 4.375 ;
        RECT  7.045 2.570 7.075 2.925 ;
        RECT  6.985 2.570 7.045 3.065 ;
        RECT  6.755 0.630 6.985 3.065 ;
        RECT  6.465 1.405 6.755 1.635 ;
        RECT  2.535 2.835 6.755 3.065 ;
        RECT  6.295 0.675 6.525 1.090 ;
        RECT  3.600 0.675 6.295 0.905 ;
        RECT  5.640 3.295 6.015 3.645 ;
        RECT  3.210 3.295 5.640 3.525 ;
        RECT  3.240 1.135 5.260 1.365 ;
        RECT  1.860 2.375 4.940 2.605 ;
        RECT  3.010 0.750 3.240 1.365 ;
        RECT  2.980 3.295 3.210 3.830 ;
        RECT  2.900 0.750 3.010 1.090 ;
        RECT  2.870 3.490 2.980 3.830 ;
        RECT  2.305 2.835 2.535 3.505 ;
        RECT  0.520 3.275 2.305 3.505 ;
        RECT  1.730 2.375 1.860 3.045 ;
        RECT  1.500 1.260 1.730 3.045 ;
        RECT  0.395 2.780 0.520 3.505 ;
        RECT  0.395 1.325 0.465 1.680 ;
        RECT  0.290 1.325 0.395 3.505 ;
        RECT  0.165 1.325 0.290 3.145 ;
    END
END EDFFTRX4

MACRO EDFFTRX2
    CLASS CORE ;
    FOREIGN EDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFTRXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 4.060 2.500 4.340 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.165 2.935 17.525 3.275 ;
        RECT  16.935 0.735 17.165 3.755 ;
        RECT  16.660 0.735 16.935 0.965 ;
        RECT  16.715 3.525 16.935 3.755 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.475 1.195 16.705 3.100 ;
        RECT  16.285 1.195 16.475 1.540 ;
        RECT  16.170 2.870 16.475 3.100 ;
        RECT  15.330 1.195 16.285 1.425 ;
        RECT  15.935 2.870 16.170 4.315 ;
        RECT  15.745 2.870 15.935 3.210 ;
        RECT  15.395 4.085 15.935 4.315 ;
        RECT  15.100 1.045 15.330 1.425 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.825 1.715 5.020 1.945 ;
        RECT  4.595 1.715 4.825 2.095 ;
        RECT  4.405 1.820 4.595 2.095 ;
        RECT  3.745 1.865 4.405 2.095 ;
        RECT  3.405 1.820 3.745 2.160 ;
        RECT  3.085 1.820 3.405 2.110 ;
        RECT  2.855 1.845 3.085 2.155 ;
        RECT  1.910 1.870 2.855 2.155 ;
        RECT  1.680 1.870 1.910 2.210 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.230 2.380 5.800 2.665 ;
        RECT  4.890 2.330 5.230 2.670 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.985 2.965 1.105 3.195 ;
        RECT  0.830 2.415 0.985 3.195 ;
        RECT  0.755 2.030 0.830 3.195 ;
        RECT  0.600 2.030 0.755 2.645 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.240 -0.400 17.820 0.400 ;
        RECT  15.900 -0.400 16.240 0.575 ;
        RECT  14.020 -0.400 15.900 0.400 ;
        RECT  13.680 -0.400 14.020 0.575 ;
        RECT  11.065 -0.400 13.680 0.400 ;
        RECT  10.835 -0.400 11.065 1.365 ;
        RECT  8.130 -0.400 10.835 0.400 ;
        RECT  7.900 -0.400 8.130 0.900 ;
        RECT  1.760 -0.400 7.900 0.400 ;
        RECT  1.420 -0.400 1.760 0.575 ;
        RECT  0.000 -0.400 1.420 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.805 4.640 17.820 5.440 ;
        RECT  16.465 4.090 16.805 5.440 ;
        RECT  14.600 4.640 16.465 5.440 ;
        RECT  14.370 3.590 14.600 5.440 ;
        RECT  12.795 4.640 14.370 5.440 ;
        RECT  12.455 4.465 12.795 5.440 ;
        RECT  10.155 4.640 12.455 5.440 ;
        RECT  9.815 4.465 10.155 5.440 ;
        RECT  7.640 4.640 9.815 5.440 ;
        RECT  7.300 4.465 7.640 5.440 ;
        RECT  4.150 4.640 7.300 5.440 ;
        RECT  3.810 4.465 4.150 5.440 ;
        RECT  1.260 4.640 3.810 5.440 ;
        RECT  0.920 4.465 1.260 5.440 ;
        RECT  0.000 4.640 0.920 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.015 1.920 16.245 2.335 ;
        RECT  15.405 2.105 16.015 2.335 ;
        RECT  15.380 1.655 15.405 3.215 ;
        RECT  15.175 1.655 15.380 3.660 ;
        RECT  14.685 1.655 15.175 1.885 ;
        RECT  15.040 2.985 15.175 3.660 ;
        RECT  14.070 2.985 15.040 3.215 ;
        RECT  14.715 2.120 14.945 2.575 ;
        RECT  12.620 2.345 14.715 2.575 ;
        RECT  14.450 1.220 14.685 1.885 ;
        RECT  14.345 1.220 14.450 1.560 ;
        RECT  13.840 2.985 14.070 4.360 ;
        RECT  12.200 3.945 13.840 4.175 ;
        RECT  12.700 3.275 13.295 3.505 ;
        RECT  11.525 0.705 13.040 0.935 ;
        RECT  12.620 3.275 12.700 3.655 ;
        RECT  12.620 1.460 12.675 1.800 ;
        RECT  12.390 1.460 12.620 3.655 ;
        RECT  12.335 1.460 12.390 1.800 ;
        RECT  11.640 3.425 12.390 3.655 ;
        RECT  11.970 3.945 12.200 4.410 ;
        RECT  10.615 4.180 11.970 4.410 ;
        RECT  11.410 3.425 11.640 3.825 ;
        RECT  11.475 0.705 11.525 2.025 ;
        RECT  11.295 0.705 11.475 2.965 ;
        RECT  11.135 3.595 11.410 3.825 ;
        RECT  11.245 1.795 11.295 2.965 ;
        RECT  11.220 2.735 11.245 2.965 ;
        RECT  10.850 2.735 11.220 3.105 ;
        RECT  10.375 2.735 10.850 2.965 ;
        RECT  10.385 4.000 10.615 4.410 ;
        RECT  10.375 0.640 10.600 1.925 ;
        RECT  3.540 4.000 10.385 4.230 ;
        RECT  10.370 0.640 10.375 2.965 ;
        RECT  8.590 0.640 10.370 0.870 ;
        RECT  10.145 1.640 10.370 2.965 ;
        RECT  9.945 2.735 10.145 2.965 ;
        RECT  9.715 1.100 10.135 1.330 ;
        RECT  9.715 2.735 9.945 3.110 ;
        RECT  9.580 1.100 9.715 2.095 ;
        RECT  9.485 1.100 9.580 2.460 ;
        RECT  9.350 1.100 9.485 3.765 ;
        RECT  9.255 2.230 9.350 3.765 ;
        RECT  9.050 3.535 9.255 3.765 ;
        RECT  8.875 1.310 9.050 2.000 ;
        RECT  8.875 2.610 9.025 2.975 ;
        RECT  8.820 1.310 8.875 3.300 ;
        RECT  8.645 1.770 8.820 3.300 ;
        RECT  8.585 1.770 8.645 2.165 ;
        RECT  8.435 3.070 8.645 3.300 ;
        RECT  8.360 0.640 8.590 1.395 ;
        RECT  7.980 1.935 8.585 2.165 ;
        RECT  8.125 3.070 8.435 3.680 ;
        RECT  8.070 2.455 8.415 2.835 ;
        RECT  7.425 1.165 8.360 1.395 ;
        RECT  8.070 3.450 8.125 3.680 ;
        RECT  7.090 2.455 8.070 2.685 ;
        RECT  7.640 1.880 7.980 2.220 ;
        RECT  7.195 0.635 7.425 1.395 ;
        RECT  6.505 0.635 7.195 0.865 ;
        RECT  6.965 2.065 7.090 3.595 ;
        RECT  6.860 1.095 6.965 3.595 ;
        RECT  6.735 1.095 6.860 2.295 ;
        RECT  5.800 3.365 6.860 3.595 ;
        RECT  6.325 2.715 6.625 3.135 ;
        RECT  6.380 0.635 6.505 1.655 ;
        RECT  6.325 0.635 6.380 1.860 ;
        RECT  6.275 0.635 6.325 3.135 ;
        RECT  6.095 1.425 6.275 3.135 ;
        RECT  6.040 1.520 6.095 1.860 ;
        RECT  2.270 2.905 6.095 3.135 ;
        RECT  5.815 0.630 6.045 1.190 ;
        RECT  3.765 0.630 5.815 0.860 ;
        RECT  2.735 3.365 5.415 3.595 ;
        RECT  4.365 1.095 4.740 1.325 ;
        RECT  4.405 2.330 4.460 2.670 ;
        RECT  4.120 2.330 4.405 2.675 ;
        RECT  4.135 1.095 4.365 1.590 ;
        RECT  2.730 1.360 4.135 1.590 ;
        RECT  1.810 2.445 4.120 2.675 ;
        RECT  3.535 0.630 3.765 1.130 ;
        RECT  3.310 4.000 3.540 4.265 ;
        RECT  3.040 0.900 3.535 1.130 ;
        RECT  2.980 4.035 3.310 4.265 ;
        RECT  2.505 3.365 2.735 3.800 ;
        RECT  2.500 0.665 2.730 1.590 ;
        RECT  2.340 0.665 2.500 0.895 ;
        RECT  2.040 2.905 2.270 3.730 ;
        RECT  0.520 3.500 2.040 3.730 ;
        RECT  1.540 1.290 1.880 1.630 ;
        RECT  1.580 2.445 1.810 3.100 ;
        RECT  1.450 2.445 1.580 2.675 ;
        RECT  1.450 1.400 1.540 1.630 ;
        RECT  1.220 1.400 1.450 2.675 ;
        RECT  0.370 1.200 0.520 1.540 ;
        RECT  0.370 2.875 0.520 3.730 ;
        RECT  0.180 1.200 0.370 3.730 ;
        RECT  0.140 1.255 0.180 3.730 ;
    END
END EDFFTRX2

MACRO EDFFTRX1
    CLASS CORE ;
    FOREIGN EDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFTRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 4.015 2.120 4.340 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.795 3.520 15.905 3.860 ;
        RECT  15.625 3.135 15.795 3.860 ;
        RECT  15.565 2.075 15.625 3.860 ;
        RECT  15.535 2.075 15.565 3.365 ;
        RECT  15.395 1.350 15.535 3.365 ;
        RECT  15.305 1.350 15.395 2.385 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.845 1.025 15.075 3.520 ;
        RECT  14.650 1.025 14.845 1.255 ;
        RECT  14.660 3.195 14.845 3.520 ;
        RECT  14.465 3.290 14.660 3.520 ;
        RECT  14.475 0.740 14.650 1.255 ;
        RECT  14.420 0.685 14.475 1.255 ;
        RECT  14.235 3.290 14.465 4.315 ;
        RECT  14.135 0.685 14.420 1.025 ;
        RECT  14.125 3.510 14.235 4.315 ;
        RECT  14.075 4.085 14.125 4.315 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 1.815 5.025 2.045 ;
        RECT  2.855 1.815 3.085 2.155 ;
        RECT  1.850 1.865 2.855 2.155 ;
        RECT  1.620 1.810 1.850 2.155 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 1.845 5.725 2.535 ;
        RECT  5.355 2.305 5.420 2.535 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 2.965 1.105 3.195 ;
        RECT  0.855 2.370 0.925 3.195 ;
        RECT  0.695 2.030 0.855 3.195 ;
        RECT  0.625 2.030 0.695 2.600 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.465 -0.400 16.500 0.400 ;
        RECT  15.125 -0.400 15.465 0.575 ;
        RECT  13.755 -0.400 15.125 0.400 ;
        RECT  13.415 -0.400 13.755 0.955 ;
        RECT  11.060 -0.400 13.415 0.400 ;
        RECT  10.830 -0.400 11.060 1.415 ;
        RECT  8.200 -0.400 10.830 0.400 ;
        RECT  7.860 -0.400 8.200 0.885 ;
        RECT  1.765 -0.400 7.860 0.400 ;
        RECT  1.425 -0.400 1.765 0.575 ;
        RECT  0.000 -0.400 1.425 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.185 4.640 16.500 5.440 ;
        RECT  14.845 3.755 15.185 5.440 ;
        RECT  12.910 4.640 14.845 5.440 ;
        RECT  12.680 3.310 12.910 5.440 ;
        RECT  10.270 4.640 12.680 5.440 ;
        RECT  9.930 4.465 10.270 5.440 ;
        RECT  7.740 4.640 9.930 5.440 ;
        RECT  7.400 4.465 7.740 5.440 ;
        RECT  4.170 4.640 7.400 5.440 ;
        RECT  3.830 4.465 4.170 5.440 ;
        RECT  1.130 4.640 3.830 5.440 ;
        RECT  0.790 4.465 1.130 5.440 ;
        RECT  0.000 4.640 0.790 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.460 2.200 14.615 2.560 ;
        RECT  14.460 1.495 14.515 1.835 ;
        RECT  14.390 1.495 14.460 2.560 ;
        RECT  14.175 1.495 14.390 3.060 ;
        RECT  14.160 1.550 14.175 3.060 ;
        RECT  13.605 2.830 14.160 3.060 ;
        RECT  13.590 2.010 13.930 2.350 ;
        RECT  13.605 3.320 13.690 3.660 ;
        RECT  13.375 2.830 13.605 3.660 ;
        RECT  13.415 2.010 13.590 2.240 ;
        RECT  13.185 1.765 13.415 2.240 ;
        RECT  12.405 2.830 13.375 3.060 ;
        RECT  13.350 3.320 13.375 3.660 ;
        RECT  12.410 1.765 13.185 1.995 ;
        RECT  11.785 0.705 12.765 0.935 ;
        RECT  12.255 1.305 12.410 1.995 ;
        RECT  12.175 2.830 12.405 4.175 ;
        RECT  12.025 1.305 12.255 2.510 ;
        RECT  2.955 3.945 12.175 4.175 ;
        RECT  11.735 2.280 12.025 2.510 ;
        RECT  11.555 0.705 11.785 2.040 ;
        RECT  11.505 2.280 11.735 3.600 ;
        RECT  10.560 1.810 11.555 2.040 ;
        RECT  11.260 3.370 11.505 3.600 ;
        RECT  10.890 2.635 11.250 3.005 ;
        RECT  10.560 2.635 10.890 2.865 ;
        RECT  10.330 0.675 10.560 2.865 ;
        RECT  8.675 0.675 10.330 0.905 ;
        RECT  10.105 1.610 10.330 1.975 ;
        RECT  10.075 2.635 10.330 2.865 ;
        RECT  9.615 1.135 10.100 1.365 ;
        RECT  9.845 2.635 10.075 3.115 ;
        RECT  9.385 1.135 9.615 3.650 ;
        RECT  9.285 1.135 9.385 1.560 ;
        RECT  9.225 3.310 9.385 3.650 ;
        RECT  8.995 2.610 9.150 2.975 ;
        RECT  8.740 1.580 9.005 1.810 ;
        RECT  8.765 2.195 8.995 3.655 ;
        RECT  8.740 2.195 8.765 2.425 ;
        RECT  7.965 3.425 8.765 3.655 ;
        RECT  8.510 1.580 8.740 2.425 ;
        RECT  8.445 0.675 8.675 1.345 ;
        RECT  7.210 2.835 8.535 3.065 ;
        RECT  7.925 2.195 8.510 2.425 ;
        RECT  7.465 1.115 8.445 1.345 ;
        RECT  7.695 2.060 7.925 2.425 ;
        RECT  7.235 0.685 7.465 1.345 ;
        RECT  6.510 0.685 7.235 0.915 ;
        RECT  6.980 2.065 7.210 3.635 ;
        RECT  6.970 2.065 6.980 2.295 ;
        RECT  5.985 3.405 6.980 3.635 ;
        RECT  6.740 1.145 6.970 2.295 ;
        RECT  6.260 2.750 6.740 3.095 ;
        RECT  6.280 0.685 6.510 1.630 ;
        RECT  6.260 1.400 6.280 1.630 ;
        RECT  6.030 1.400 6.260 3.095 ;
        RECT  5.820 0.815 6.050 1.155 ;
        RECT  5.115 2.765 6.030 2.995 ;
        RECT  3.045 0.815 5.820 1.045 ;
        RECT  2.710 3.445 5.440 3.675 ;
        RECT  4.885 2.765 5.115 3.215 ;
        RECT  2.245 2.985 4.885 3.215 ;
        RECT  2.805 1.275 4.745 1.505 ;
        RECT  1.785 2.520 4.320 2.750 ;
        RECT  2.575 0.665 2.805 1.505 ;
        RECT  2.480 3.445 2.710 3.860 ;
        RECT  2.345 0.665 2.575 0.895 ;
        RECT  2.015 2.985 2.245 3.690 ;
        RECT  0.465 3.460 2.015 3.690 ;
        RECT  1.390 1.275 1.885 1.505 ;
        RECT  1.555 2.385 1.785 3.100 ;
        RECT  1.390 2.385 1.555 2.615 ;
        RECT  1.160 1.275 1.390 2.615 ;
        RECT  0.395 1.200 0.520 1.540 ;
        RECT  0.395 2.855 0.465 3.690 ;
        RECT  0.235 1.200 0.395 3.690 ;
        RECT  0.180 1.200 0.235 3.170 ;
        RECT  0.165 1.255 0.180 3.170 ;
    END
END EDFFTRX1

MACRO EDFFXL
    CLASS CORE ;
    FOREIGN EDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.940 1.845 14.965 2.075 ;
        RECT  14.750 1.355 14.940 2.845 ;
        RECT  14.710 1.280 14.750 2.845 ;
        RECT  14.660 1.280 14.710 1.820 ;
        RECT  14.550 2.615 14.710 2.845 ;
        RECT  14.410 1.280 14.660 1.620 ;
        RECT  14.320 2.615 14.550 3.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.825 0.885 14.055 3.755 ;
        RECT  13.245 0.885 13.825 1.115 ;
        RECT  13.720 3.500 13.825 3.755 ;
        RECT  13.565 3.525 13.720 3.755 ;
        RECT  13.335 3.525 13.565 4.145 ;
        RECT  12.765 3.915 13.335 4.145 ;
        RECT  13.015 0.725 13.245 1.115 ;
        RECT  12.495 0.725 13.015 0.955 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 3.970 2.090 4.380 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.975 2.405 5.065 2.635 ;
        RECT  4.745 2.145 4.975 2.635 ;
        RECT  4.540 2.145 4.745 2.375 ;
        RECT  4.310 1.980 4.540 2.375 ;
        RECT  4.110 1.980 4.310 2.210 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.885 2.380 1.175 2.660 ;
        RECT  0.655 2.120 0.885 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.985 -0.400 15.180 0.400 ;
        RECT  13.645 -0.400 13.985 0.575 ;
        RECT  12.030 -0.400 13.645 0.400 ;
        RECT  11.690 -0.400 12.030 0.575 ;
        RECT  9.350 -0.400 11.690 0.400 ;
        RECT  9.010 -0.400 9.350 1.060 ;
        RECT  7.050 -0.400 9.010 0.400 ;
        RECT  6.710 -0.400 7.050 1.240 ;
        RECT  3.530 -0.400 6.710 0.400 ;
        RECT  3.190 -0.400 3.530 0.575 ;
        RECT  0.890 -0.400 3.190 0.400 ;
        RECT  0.550 -0.400 0.890 0.575 ;
        RECT  0.000 -0.400 0.550 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.890 4.640 15.180 5.440 ;
        RECT  13.550 4.465 13.890 5.440 ;
        RECT  12.335 4.640 13.550 5.440 ;
        RECT  11.995 4.465 12.335 5.440 ;
        RECT  8.895 4.640 11.995 5.440 ;
        RECT  8.555 4.465 8.895 5.440 ;
        RECT  7.495 4.640 8.555 5.440 ;
        RECT  7.155 4.465 7.495 5.440 ;
        RECT  4.100 4.640 7.155 5.440 ;
        RECT  3.760 4.465 4.100 5.440 ;
        RECT  1.120 4.640 3.760 5.440 ;
        RECT  0.780 4.465 1.120 5.440 ;
        RECT  0.000 4.640 0.780 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.305 1.490 13.535 3.260 ;
        RECT  12.535 1.490 13.305 1.720 ;
        RECT  11.825 3.030 13.305 3.260 ;
        RECT  10.835 2.095 12.485 2.325 ;
        RECT  11.750 3.030 11.825 4.225 ;
        RECT  11.595 3.030 11.750 4.310 ;
        RECT  11.520 3.995 11.595 4.310 ;
        RECT  2.525 3.995 11.520 4.225 ;
        RECT  9.945 0.685 11.030 0.915 ;
        RECT  10.615 2.095 10.835 3.730 ;
        RECT  10.605 1.330 10.615 3.730 ;
        RECT  10.385 1.330 10.605 2.325 ;
        RECT  10.455 3.500 10.605 3.730 ;
        RECT  9.945 2.610 10.370 2.960 ;
        RECT  9.715 0.685 9.945 3.670 ;
        RECT  5.660 3.440 9.715 3.670 ;
        RECT  9.250 1.310 9.480 3.135 ;
        RECT  8.495 1.310 9.250 1.540 ;
        RECT  8.555 2.905 9.250 3.135 ;
        RECT  8.065 2.335 9.015 2.565 ;
        RECT  8.265 0.655 8.495 1.540 ;
        RECT  8.055 0.655 8.265 0.885 ;
        RECT  8.050 2.335 8.065 3.065 ;
        RECT  7.820 1.775 8.050 3.065 ;
        RECT  7.795 1.775 7.820 2.005 ;
        RECT  7.715 2.835 7.820 3.065 ;
        RECT  7.565 0.900 7.795 2.005 ;
        RECT  7.360 2.235 7.590 2.590 ;
        RECT  6.590 1.555 7.565 1.785 ;
        RECT  6.120 2.235 7.360 2.465 ;
        RECT  6.360 1.555 6.590 1.920 ;
        RECT  5.890 1.025 6.120 3.110 ;
        RECT  5.690 1.025 5.890 1.255 ;
        RECT  5.350 0.915 5.690 1.255 ;
        RECT  5.430 1.520 5.660 3.670 ;
        RECT  4.075 1.520 5.430 1.750 ;
        RECT  4.970 2.895 5.200 3.715 ;
        RECT  2.245 3.405 4.970 3.635 ;
        RECT  4.655 0.970 4.890 1.200 ;
        RECT  4.425 0.805 4.655 1.200 ;
        RECT  2.455 0.805 4.425 1.035 ;
        RECT  3.155 2.685 4.175 2.915 ;
        RECT  3.845 1.270 4.075 1.750 ;
        RECT  0.520 1.270 3.845 1.500 ;
        RECT  2.925 2.050 3.155 2.915 ;
        RECT  1.985 2.050 2.925 2.280 ;
        RECT  2.225 0.795 2.455 1.035 ;
        RECT  1.820 0.795 2.225 1.025 ;
        RECT  1.955 1.735 1.985 2.280 ;
        RECT  1.725 1.735 1.955 3.575 ;
        RECT  1.580 1.735 1.725 1.965 ;
        RECT  1.540 3.345 1.725 3.575 ;
        RECT  0.405 1.270 0.520 1.660 ;
        RECT  0.405 3.475 0.520 3.705 ;
        RECT  0.235 1.270 0.405 3.705 ;
        RECT  0.180 1.320 0.235 3.705 ;
        RECT  0.175 1.375 0.180 3.705 ;
    END
END EDFFXL

MACRO EDFFX4
    CLASS CORE ;
    FOREIGN EDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.000 1.460 19.585 1.800 ;
        RECT  19.000 2.900 19.505 3.240 ;
        RECT  18.620 1.260 19.000 3.240 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.960 1.260 18.340 3.240 ;
        RECT  17.885 2.900 17.960 3.240 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 1.420 3.745 2.075 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.865 2.405 5.065 2.635 ;
        RECT  4.635 1.620 4.865 2.635 ;
        RECT  4.395 1.620 4.635 1.850 ;
        RECT  4.055 1.510 4.395 1.850 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.025 0.520 2.655 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.225 -0.400 20.460 0.400 ;
        RECT  19.885 -0.400 20.225 1.050 ;
        RECT  18.945 -0.400 19.885 0.400 ;
        RECT  18.605 -0.400 18.945 0.995 ;
        RECT  17.665 -0.400 18.605 0.400 ;
        RECT  17.325 -0.400 17.665 1.050 ;
        RECT  16.240 -0.400 17.325 0.400 ;
        RECT  15.900 -0.400 16.240 1.625 ;
        RECT  13.130 -0.400 15.900 0.400 ;
        RECT  12.790 -0.400 13.130 0.575 ;
        RECT  10.290 -0.400 12.790 0.400 ;
        RECT  9.950 -0.400 10.290 0.575 ;
        RECT  8.460 -0.400 9.950 0.400 ;
        RECT  8.230 -0.400 8.460 1.300 ;
        RECT  6.950 -0.400 8.230 0.400 ;
        RECT  6.610 -0.400 6.950 1.155 ;
        RECT  3.410 -0.400 6.610 0.400 ;
        RECT  3.070 -0.400 3.410 0.575 ;
        RECT  1.240 -0.400 3.070 0.400 ;
        RECT  0.900 -0.400 1.240 0.950 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.145 4.640 20.460 5.440 ;
        RECT  19.805 4.090 20.145 5.440 ;
        RECT  18.865 4.640 19.805 5.440 ;
        RECT  18.525 4.090 18.865 5.440 ;
        RECT  17.235 4.640 18.525 5.440 ;
        RECT  16.895 4.090 17.235 5.440 ;
        RECT  15.585 4.640 16.895 5.440 ;
        RECT  15.245 4.465 15.585 5.440 ;
        RECT  12.805 4.640 15.245 5.440 ;
        RECT  12.465 4.465 12.805 5.440 ;
        RECT  10.000 4.640 12.465 5.440 ;
        RECT  9.660 4.465 10.000 5.440 ;
        RECT  7.570 4.640 9.660 5.440 ;
        RECT  7.230 4.465 7.570 5.440 ;
        RECT  4.065 4.640 7.230 5.440 ;
        RECT  3.725 4.465 4.065 5.440 ;
        RECT  1.410 4.640 3.725 5.440 ;
        RECT  1.070 4.465 1.410 5.440 ;
        RECT  0.000 4.640 1.070 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.735 2.440 19.965 3.805 ;
        RECT  19.665 2.440 19.735 2.670 ;
        RECT  17.645 3.575 19.735 3.805 ;
        RECT  19.435 2.055 19.665 2.670 ;
        RECT  17.415 1.460 17.645 3.805 ;
        RECT  16.910 1.460 17.415 1.690 ;
        RECT  16.500 3.575 17.415 3.805 ;
        RECT  15.265 2.035 17.120 2.265 ;
        RECT  16.680 0.870 16.910 1.690 ;
        RECT  16.270 3.575 16.500 4.085 ;
        RECT  15.725 3.855 16.270 4.085 ;
        RECT  15.495 2.620 15.725 4.235 ;
        RECT  2.440 4.005 15.495 4.235 ;
        RECT  15.035 1.265 15.265 3.655 ;
        RECT  14.505 1.265 15.035 1.495 ;
        RECT  11.430 3.425 15.035 3.655 ;
        RECT  14.575 2.085 14.805 3.135 ;
        RECT  13.705 2.905 14.575 3.135 ;
        RECT  14.275 0.865 14.505 1.495 ;
        RECT  11.470 0.865 14.275 1.095 ;
        RECT  13.055 1.740 14.085 1.970 ;
        RECT  13.475 2.540 13.705 3.135 ;
        RECT  12.415 2.905 13.475 3.135 ;
        RECT  12.825 1.735 13.055 1.970 ;
        RECT  10.465 1.735 12.825 1.965 ;
        RECT  12.185 2.745 12.415 3.135 ;
        RECT  11.025 2.745 12.185 2.975 ;
        RECT  11.200 3.290 11.430 3.655 ;
        RECT  10.930 2.535 11.025 2.975 ;
        RECT  10.700 2.535 10.930 3.655 ;
        RECT  8.575 3.425 10.700 3.655 ;
        RECT  10.235 1.335 10.465 3.075 ;
        RECT  10.225 1.335 10.235 1.965 ;
        RECT  8.720 2.845 10.235 3.075 ;
        RECT  9.530 1.335 10.225 1.565 ;
        RECT  9.775 2.220 10.005 2.615 ;
        RECT  8.350 2.385 9.775 2.615 ;
        RECT  9.475 1.255 9.530 1.565 ;
        RECT  9.245 0.630 9.475 1.565 ;
        RECT  8.720 0.630 9.245 0.860 ;
        RECT  8.345 3.425 8.575 3.770 ;
        RECT  8.295 2.385 8.350 3.075 ;
        RECT  5.895 3.540 8.345 3.770 ;
        RECT  8.185 2.320 8.295 3.075 ;
        RECT  7.995 2.275 8.185 3.075 ;
        RECT  7.965 2.275 7.995 2.550 ;
        RECT  7.735 0.925 7.965 2.550 ;
        RECT  7.410 0.925 7.735 1.155 ;
        RECT  7.380 2.320 7.735 2.550 ;
        RECT  6.415 1.465 7.425 1.695 ;
        RECT  7.040 2.210 7.380 2.550 ;
        RECT  6.355 1.465 6.415 3.110 ;
        RECT  6.185 0.760 6.355 3.110 ;
        RECT  6.125 0.760 6.185 1.700 ;
        RECT  5.110 0.760 6.125 0.990 ;
        RECT  5.665 1.745 5.895 3.770 ;
        RECT  5.100 1.745 5.665 1.975 ;
        RECT  0.980 3.540 5.665 3.770 ;
        RECT  5.080 2.965 5.310 3.305 ;
        RECT  2.485 3.075 5.080 3.305 ;
        RECT  4.390 0.660 4.730 1.040 ;
        RECT  2.455 0.810 4.390 1.040 ;
        RECT  4.285 2.285 4.350 2.570 ;
        RECT  4.000 2.285 4.285 2.615 ;
        RECT  2.975 2.385 4.000 2.615 ;
        RECT  2.745 1.405 2.975 2.615 ;
        RECT  2.510 1.405 2.745 1.735 ;
        RECT  1.695 1.505 2.510 1.735 ;
        RECT  2.255 2.850 2.485 3.305 ;
        RECT  2.225 0.730 2.455 1.040 ;
        RECT  1.600 0.730 2.225 0.960 ;
        RECT  1.695 2.835 1.840 3.065 ;
        RECT  1.465 1.505 1.695 3.065 ;
        RECT  0.750 1.400 0.980 3.770 ;
        RECT  0.520 1.400 0.750 1.630 ;
        RECT  0.520 2.890 0.750 3.770 ;
        RECT  0.180 0.820 0.520 1.630 ;
        RECT  0.180 2.890 0.520 4.170 ;
    END
END EDFFX4

MACRO EDFFX2
    CLASS CORE ;
    FOREIGN EDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.320 1.340 17.375 1.680 ;
        RECT  17.090 1.340 17.320 3.095 ;
        RECT  17.035 1.340 17.090 1.680 ;
        RECT  17.015 2.755 17.090 3.095 ;
        RECT  16.865 2.755 17.015 3.755 ;
        RECT  16.785 2.810 16.865 3.755 ;
        RECT  16.715 3.525 16.785 3.755 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.980 2.965 16.285 3.195 ;
        RECT  15.840 2.940 15.980 3.195 ;
        RECT  15.705 1.445 15.900 1.675 ;
        RECT  15.705 2.755 15.840 3.195 ;
        RECT  15.475 1.445 15.705 3.195 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 3.950 2.000 4.380 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.975 2.405 5.065 2.635 ;
        RECT  4.745 2.145 4.975 2.635 ;
        RECT  4.235 2.145 4.745 2.375 ;
        RECT  4.005 2.055 4.235 2.375 ;
        RECT  3.885 2.055 4.005 2.285 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.120 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.610 -0.400 17.820 0.400 ;
        RECT  16.270 -0.400 16.610 0.575 ;
        RECT  14.400 -0.400 16.270 0.400 ;
        RECT  14.060 -0.400 14.400 0.575 ;
        RECT  12.815 -0.400 14.060 0.400 ;
        RECT  12.475 -0.400 12.815 0.575 ;
        RECT  10.010 -0.400 12.475 0.400 ;
        RECT  9.670 -0.400 10.010 1.295 ;
        RECT  6.915 -0.400 9.670 0.400 ;
        RECT  6.575 -0.400 6.915 1.300 ;
        RECT  3.385 -0.400 6.575 0.400 ;
        RECT  3.045 -0.400 3.385 0.575 ;
        RECT  0.760 -0.400 3.045 0.400 ;
        RECT  0.420 -0.400 0.760 0.575 ;
        RECT  0.000 -0.400 0.420 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.525 4.640 17.820 5.440 ;
        RECT  16.185 4.465 16.525 5.440 ;
        RECT  14.080 4.640 16.185 5.440 ;
        RECT  13.740 4.465 14.080 5.440 ;
        RECT  12.830 4.640 13.740 5.440 ;
        RECT  12.490 4.465 12.830 5.440 ;
        RECT  9.220 4.640 12.490 5.440 ;
        RECT  8.880 4.465 9.220 5.440 ;
        RECT  7.545 4.640 8.880 5.440 ;
        RECT  7.205 4.465 7.545 5.440 ;
        RECT  3.985 4.640 7.205 5.440 ;
        RECT  3.645 4.465 3.985 5.440 ;
        RECT  1.065 4.640 3.645 5.440 ;
        RECT  1.065 3.335 1.240 3.565 ;
        RECT  0.835 3.335 1.065 5.440 ;
        RECT  0.000 4.640 0.835 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.585 1.915 16.815 2.280 ;
        RECT  16.415 1.915 16.585 2.145 ;
        RECT  16.185 0.915 16.415 2.145 ;
        RECT  15.200 0.915 16.185 1.145 ;
        RECT  15.115 0.685 15.200 1.145 ;
        RECT  15.065 0.685 15.115 3.290 ;
        RECT  14.885 0.685 15.065 4.175 ;
        RECT  14.855 0.685 14.885 1.145 ;
        RECT  14.835 3.060 14.885 4.175 ;
        RECT  2.565 3.945 14.835 4.175 ;
        RECT  13.675 2.220 14.650 2.575 ;
        RECT  13.445 1.265 13.675 3.325 ;
        RECT  12.830 1.265 13.445 1.495 ;
        RECT  11.360 3.095 13.445 3.325 ;
        RECT  12.985 1.790 13.215 2.785 ;
        RECT  10.585 2.555 12.985 2.785 ;
        RECT  12.600 1.245 12.830 1.495 ;
        RECT  10.950 1.245 12.600 1.475 ;
        RECT  11.130 3.095 11.360 3.575 ;
        RECT  9.995 1.835 11.280 2.065 ;
        RECT  10.955 3.345 11.130 3.575 ;
        RECT  10.355 2.555 10.585 3.705 ;
        RECT  6.495 3.475 10.355 3.705 ;
        RECT  9.985 1.695 9.995 2.065 ;
        RECT  9.755 1.695 9.985 3.245 ;
        RECT  8.910 1.695 9.755 1.925 ;
        RECT  8.940 3.015 9.755 3.245 ;
        RECT  8.325 2.305 9.265 2.535 ;
        RECT  8.680 0.675 8.910 1.925 ;
        RECT  8.070 0.675 8.680 0.905 ;
        RECT  8.195 2.305 8.325 3.075 ;
        RECT  7.965 1.825 8.195 3.075 ;
        RECT  7.585 1.825 7.965 2.055 ;
        RECT  6.170 2.295 7.700 2.525 ;
        RECT  7.355 0.965 7.585 2.055 ;
        RECT  6.635 1.825 7.355 2.055 ;
        RECT  6.405 1.680 6.635 2.055 ;
        RECT  6.180 3.425 6.495 3.705 ;
        RECT  5.710 3.425 6.180 3.655 ;
        RECT  5.940 0.905 6.170 3.110 ;
        RECT  5.260 0.905 5.940 1.235 ;
        RECT  5.480 1.605 5.710 3.655 ;
        RECT  4.775 1.605 5.480 1.835 ;
        RECT  5.205 0.905 5.260 1.135 ;
        RECT  5.020 3.265 5.250 3.650 ;
        RECT  4.610 3.265 5.020 3.575 ;
        RECT  4.545 1.265 4.775 1.835 ;
        RECT  2.815 0.805 4.745 1.035 ;
        RECT  2.325 3.345 4.610 3.575 ;
        RECT  2.355 1.265 4.545 1.495 ;
        RECT  3.155 2.775 4.265 3.005 ;
        RECT  2.925 2.145 3.155 3.005 ;
        RECT  1.910 2.145 2.925 2.375 ;
        RECT  2.585 0.735 2.815 1.035 ;
        RECT  1.680 0.735 2.585 0.965 ;
        RECT  2.125 1.195 2.355 1.495 ;
        RECT  0.520 1.195 2.125 1.425 ;
        RECT  1.680 1.655 1.910 3.620 ;
        RECT  1.665 1.655 1.680 2.375 ;
        RECT  1.540 1.655 1.665 1.885 ;
        RECT  0.405 1.195 0.520 1.660 ;
        RECT  0.405 3.425 0.520 3.655 ;
        RECT  0.235 1.195 0.405 3.655 ;
        RECT  0.180 1.320 0.235 3.655 ;
        RECT  0.175 1.375 0.180 3.655 ;
    END
END EDFFX2

MACRO EDFFX1
    CLASS CORE ;
    FOREIGN EDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.890 1.845 14.965 2.075 ;
        RECT  14.750 1.380 14.890 2.845 ;
        RECT  14.660 1.270 14.750 2.845 ;
        RECT  14.410 1.270 14.660 1.610 ;
        RECT  14.550 2.615 14.660 2.845 ;
        RECT  14.320 2.615 14.550 3.705 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.825 0.885 14.055 3.755 ;
        RECT  13.245 0.885 13.825 1.115 ;
        RECT  13.720 3.500 13.825 3.755 ;
        RECT  13.565 3.525 13.720 3.755 ;
        RECT  13.335 3.525 13.565 4.145 ;
        RECT  12.765 3.915 13.335 4.145 ;
        RECT  13.015 0.695 13.245 1.115 ;
        RECT  12.985 0.695 13.015 0.955 ;
        RECT  12.495 0.695 12.985 0.925 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 3.970 2.090 4.380 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.975 2.405 5.065 2.635 ;
        RECT  4.745 2.145 4.975 2.635 ;
        RECT  4.110 2.145 4.745 2.375 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.885 2.380 1.175 2.660 ;
        RECT  0.655 2.120 0.885 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.985 -0.400 15.180 0.400 ;
        RECT  13.645 -0.400 13.985 0.575 ;
        RECT  12.030 -0.400 13.645 0.400 ;
        RECT  11.690 -0.400 12.030 0.575 ;
        RECT  9.375 -0.400 11.690 0.400 ;
        RECT  9.035 -0.400 9.375 1.235 ;
        RECT  7.050 -0.400 9.035 0.400 ;
        RECT  6.710 -0.400 7.050 1.240 ;
        RECT  3.530 -0.400 6.710 0.400 ;
        RECT  3.190 -0.400 3.530 0.575 ;
        RECT  0.890 -0.400 3.190 0.400 ;
        RECT  0.550 -0.400 0.890 0.575 ;
        RECT  0.000 -0.400 0.550 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.890 4.640 15.180 5.440 ;
        RECT  13.550 4.465 13.890 5.440 ;
        RECT  12.335 4.640 13.550 5.440 ;
        RECT  11.995 4.465 12.335 5.440 ;
        RECT  8.895 4.640 11.995 5.440 ;
        RECT  8.555 4.465 8.895 5.440 ;
        RECT  7.495 4.640 8.555 5.440 ;
        RECT  7.155 4.465 7.495 5.440 ;
        RECT  4.100 4.640 7.155 5.440 ;
        RECT  3.760 4.465 4.100 5.440 ;
        RECT  1.120 4.640 3.760 5.440 ;
        RECT  0.780 4.465 1.120 5.440 ;
        RECT  0.000 4.640 0.780 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.305 1.490 13.535 3.255 ;
        RECT  12.535 1.490 13.305 1.720 ;
        RECT  11.825 3.025 13.305 3.255 ;
        RECT  10.835 2.095 12.485 2.325 ;
        RECT  11.750 3.025 11.825 4.225 ;
        RECT  11.595 3.025 11.750 4.310 ;
        RECT  11.520 3.995 11.595 4.310 ;
        RECT  2.525 3.995 11.520 4.225 ;
        RECT  9.945 0.685 11.030 0.915 ;
        RECT  10.605 2.095 10.835 3.575 ;
        RECT  10.600 2.095 10.605 2.325 ;
        RECT  10.455 3.345 10.605 3.575 ;
        RECT  10.370 1.330 10.600 2.325 ;
        RECT  9.945 2.610 10.370 2.960 ;
        RECT  9.715 0.685 9.945 3.670 ;
        RECT  5.660 3.440 9.715 3.670 ;
        RECT  9.250 1.470 9.480 3.135 ;
        RECT  8.520 1.470 9.250 1.700 ;
        RECT  8.525 2.905 9.250 3.135 ;
        RECT  8.065 2.335 9.015 2.565 ;
        RECT  8.290 0.675 8.520 1.700 ;
        RECT  8.055 0.675 8.290 0.905 ;
        RECT  8.050 2.335 8.065 3.055 ;
        RECT  7.820 1.555 8.050 3.055 ;
        RECT  7.795 1.555 7.820 1.785 ;
        RECT  7.715 2.825 7.820 3.055 ;
        RECT  7.565 0.900 7.795 1.785 ;
        RECT  7.360 2.235 7.590 2.590 ;
        RECT  6.590 1.555 7.565 1.785 ;
        RECT  6.120 2.235 7.360 2.465 ;
        RECT  6.360 1.555 6.590 1.920 ;
        RECT  5.890 1.025 6.120 3.110 ;
        RECT  5.690 1.025 5.890 1.255 ;
        RECT  5.350 0.915 5.690 1.255 ;
        RECT  5.430 1.625 5.660 3.670 ;
        RECT  4.075 1.625 5.430 1.855 ;
        RECT  4.970 3.230 5.200 3.635 ;
        RECT  2.245 3.405 4.970 3.635 ;
        RECT  4.655 0.970 4.890 1.200 ;
        RECT  4.425 0.805 4.655 1.200 ;
        RECT  2.455 0.805 4.425 1.035 ;
        RECT  3.155 2.855 4.175 3.085 ;
        RECT  3.845 1.270 4.075 1.855 ;
        RECT  0.520 1.270 3.845 1.500 ;
        RECT  2.925 2.145 3.155 3.085 ;
        RECT  1.955 2.145 2.925 2.375 ;
        RECT  2.225 0.725 2.455 1.035 ;
        RECT  1.820 0.725 2.225 0.955 ;
        RECT  1.890 2.145 1.955 3.575 ;
        RECT  1.725 1.735 1.890 3.575 ;
        RECT  1.605 1.735 1.725 2.375 ;
        RECT  1.540 3.345 1.725 3.575 ;
        RECT  1.550 1.735 1.605 1.965 ;
        RECT  0.405 1.270 0.520 1.660 ;
        RECT  0.405 3.425 0.520 3.655 ;
        RECT  0.235 1.270 0.405 3.655 ;
        RECT  0.180 1.320 0.235 3.655 ;
        RECT  0.175 1.375 0.180 3.655 ;
    END
END EDFFX1

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.210 1.310 4.440 3.440 ;
        RECT  4.100 1.310 4.210 1.650 ;
        RECT  4.175 2.965 4.210 3.440 ;
        RECT  4.100 3.100 4.175 3.440 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.525 1.105 3.895 ;
        RECT  0.800 3.610 0.875 3.895 ;
        RECT  0.460 3.610 0.800 3.950 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 -0.400 4.620 0.400 ;
        RECT  3.540 -0.400 3.880 0.575 ;
        RECT  1.440 -0.400 3.540 0.400 ;
        RECT  1.100 -0.400 1.440 0.575 ;
        RECT  0.000 -0.400 1.100 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 4.640 4.620 5.440 ;
        RECT  3.540 4.465 3.880 5.440 ;
        RECT  1.200 4.640 3.540 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.520 2.040 3.975 2.380 ;
        RECT  3.290 0.825 3.520 3.760 ;
        RECT  2.540 0.825 3.290 1.055 ;
        RECT  2.430 3.530 3.290 3.760 ;
        RECT  2.540 2.040 3.060 2.380 ;
        RECT  2.200 0.715 2.540 1.055 ;
        RECT  2.310 1.410 2.540 3.080 ;
        RECT  2.090 3.530 2.430 3.870 ;
        RECT  2.200 1.410 2.310 1.750 ;
        RECT  2.200 2.740 2.310 3.080 ;
        RECT  0.520 2.170 1.720 2.510 ;
        RECT  0.290 1.410 0.520 3.080 ;
        RECT  0.180 1.410 0.290 1.750 ;
        RECT  0.180 2.740 0.290 3.080 ;
    END
END DLY4X1

MACRO DLY3X1
    CLASS CORE ;
    FOREIGN DLY3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.210 1.310 4.440 3.440 ;
        RECT  4.100 1.310 4.210 1.650 ;
        RECT  4.175 2.965 4.210 3.440 ;
        RECT  4.100 3.100 4.175 3.440 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.525 1.105 3.895 ;
        RECT  0.800 3.610 0.875 3.895 ;
        RECT  0.460 3.610 0.800 3.950 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 -0.400 4.620 0.400 ;
        RECT  3.330 -0.400 3.670 0.575 ;
        RECT  1.260 -0.400 3.330 0.400 ;
        RECT  0.920 -0.400 1.260 0.575 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.680 4.640 4.620 5.440 ;
        RECT  3.330 4.465 3.680 5.440 ;
        RECT  1.260 4.640 3.330 5.440 ;
        RECT  0.920 4.465 1.260 5.440 ;
        RECT  0.000 4.640 0.920 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.410 2.040 3.955 2.380 ;
        RECT  3.180 0.825 3.410 3.760 ;
        RECT  2.430 0.825 3.180 1.055 ;
        RECT  2.430 3.530 3.180 3.760 ;
        RECT  2.420 2.040 2.950 2.380 ;
        RECT  2.090 0.715 2.430 1.055 ;
        RECT  2.090 3.530 2.430 3.870 ;
        RECT  2.190 1.410 2.420 3.080 ;
        RECT  2.080 1.410 2.190 1.750 ;
        RECT  2.080 2.740 2.190 3.080 ;
        RECT  0.520 2.170 1.780 2.510 ;
        RECT  0.290 1.410 0.520 3.080 ;
        RECT  0.180 1.410 0.290 1.750 ;
        RECT  0.180 2.740 0.290 3.080 ;
    END
END DLY3X1

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 1.310 3.780 3.440 ;
        RECT  3.440 1.310 3.550 1.650 ;
        RECT  3.515 2.965 3.550 3.440 ;
        RECT  3.440 3.100 3.515 3.440 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.525 1.105 3.895 ;
        RECT  0.800 3.610 0.875 3.895 ;
        RECT  0.460 3.610 0.800 3.950 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 -0.400 3.960 0.400 ;
        RECT  2.880 -0.400 3.220 0.575 ;
        RECT  1.260 -0.400 2.880 0.400 ;
        RECT  0.920 -0.400 1.260 0.575 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 4.640 3.960 5.440 ;
        RECT  2.880 4.465 3.220 5.440 ;
        RECT  1.260 4.640 2.880 5.440 ;
        RECT  0.920 4.465 1.260 5.440 ;
        RECT  0.000 4.640 0.920 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.210 2.040 3.315 2.380 ;
        RECT  2.980 0.825 3.210 3.760 ;
        RECT  2.240 0.825 2.980 1.055 ;
        RECT  2.240 3.530 2.980 3.760 ;
        RECT  2.240 2.040 2.700 2.380 ;
        RECT  1.900 0.715 2.240 1.055 ;
        RECT  2.010 1.410 2.240 3.080 ;
        RECT  1.900 3.530 2.240 3.870 ;
        RECT  1.900 1.410 2.010 1.750 ;
        RECT  1.900 2.740 2.010 3.080 ;
        RECT  0.520 2.170 1.720 2.510 ;
        RECT  0.290 1.410 0.520 3.080 ;
        RECT  0.180 1.410 0.290 1.750 ;
        RECT  0.180 2.740 0.290 3.080 ;
    END
END DLY2X1

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.020 3.780 1.360 ;
        RECT  3.745 3.190 3.780 3.600 ;
        RECT  3.515 1.020 3.745 3.600 ;
        RECT  3.440 1.020 3.515 1.360 ;
        RECT  3.440 3.190 3.515 3.600 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 3.500 1.180 3.780 ;
        RECT  0.790 3.470 0.875 3.780 ;
        RECT  0.450 3.470 0.790 3.810 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 -0.400 3.960 0.400 ;
        RECT  2.680 -0.400 3.020 0.575 ;
        RECT  1.420 -0.400 2.680 0.400 ;
        RECT  1.080 -0.400 1.420 0.575 ;
        RECT  0.000 -0.400 1.080 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 4.640 3.960 5.440 ;
        RECT  2.680 4.465 3.020 5.440 ;
        RECT  1.420 4.640 2.680 5.440 ;
        RECT  1.080 4.465 1.420 5.440 ;
        RECT  0.000 4.640 1.080 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.960 2.040 3.210 2.380 ;
        RECT  2.730 0.805 2.960 3.760 ;
        RECT  2.220 0.805 2.730 1.035 ;
        RECT  2.220 3.530 2.730 3.760 ;
        RECT  2.220 2.040 2.500 2.380 ;
        RECT  1.880 0.715 2.220 1.035 ;
        RECT  1.990 1.410 2.220 3.080 ;
        RECT  1.880 3.530 2.220 3.870 ;
        RECT  1.880 1.410 1.990 1.750 ;
        RECT  1.880 2.740 1.990 3.080 ;
        RECT  0.520 2.170 1.700 2.510 ;
        RECT  0.290 1.410 0.520 3.080 ;
        RECT  0.180 1.410 0.290 1.750 ;
        RECT  0.180 2.740 0.290 3.080 ;
    END
END DLY1X1

MACRO DFFTRXL
    CLASS CORE ;
    FOREIGN DFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 1.285 1.765 1.515 ;
        RECT  1.275 1.285 1.505 2.050 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.905 1.845 11.005 2.075 ;
        RECT  10.810 1.200 10.905 2.075 ;
        RECT  10.675 1.200 10.810 3.230 ;
        RECT  10.580 1.845 10.675 3.230 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 0.810 10.345 3.800 ;
        RECT  9.455 0.810 10.115 1.040 ;
        RECT  9.445 3.570 10.115 3.800 ;
        RECT  9.405 0.725 9.455 1.040 ;
        RECT  9.105 3.570 9.445 3.910 ;
        RECT  9.175 0.700 9.405 1.040 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.300 1.820 2.500 2.100 ;
        RECT  2.070 1.820 2.300 2.250 ;
        RECT  1.780 1.820 2.070 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 2.790 1.230 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.200 -0.400 11.220 0.400 ;
        RECT  9.860 -0.400 10.200 0.575 ;
        RECT  8.740 -0.400 9.860 0.400 ;
        RECT  8.400 -0.400 8.740 1.040 ;
        RECT  6.005 -0.400 8.400 0.400 ;
        RECT  5.775 -0.400 6.005 0.900 ;
        RECT  4.145 -0.400 5.775 0.400 ;
        RECT  3.915 -0.400 4.145 0.870 ;
        RECT  1.120 -0.400 3.915 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.145 4.640 11.220 5.440 ;
        RECT  10.090 4.465 10.145 5.440 ;
        RECT  9.860 4.410 10.090 5.440 ;
        RECT  9.805 4.465 9.860 5.440 ;
        RECT  8.685 4.640 9.805 5.440 ;
        RECT  8.345 3.960 8.685 5.440 ;
        RECT  6.365 4.640 8.345 5.440 ;
        RECT  6.025 3.540 6.365 5.440 ;
        RECT  4.620 4.640 6.025 5.440 ;
        RECT  4.565 4.465 4.620 5.440 ;
        RECT  4.335 4.410 4.565 5.440 ;
        RECT  4.280 4.465 4.335 5.440 ;
        RECT  1.290 4.640 4.280 5.440 ;
        RECT  0.950 4.465 1.290 5.440 ;
        RECT  0.000 4.640 0.950 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.545 1.460 9.885 3.140 ;
        RECT  9.160 1.460 9.545 1.800 ;
        RECT  9.105 2.800 9.545 3.140 ;
        RECT  8.275 1.570 9.160 1.800 ;
        RECT  8.870 2.140 9.090 2.480 ;
        RECT  8.750 2.140 8.870 2.725 ;
        RECT  8.640 2.250 8.750 2.725 ;
        RECT  7.670 2.495 8.640 2.725 ;
        RECT  8.045 1.570 8.275 2.220 ;
        RECT  7.670 3.600 7.725 3.940 ;
        RECT  7.440 1.215 7.670 3.940 ;
        RECT  7.325 1.215 7.440 1.445 ;
        RECT  7.385 3.600 7.440 3.940 ;
        RECT  7.095 1.090 7.325 1.445 ;
        RECT  6.825 1.885 7.100 2.115 ;
        RECT  6.595 1.295 6.825 3.005 ;
        RECT  5.405 1.295 6.595 1.525 ;
        RECT  5.810 2.775 6.595 3.005 ;
        RECT  5.145 1.965 6.365 2.345 ;
        RECT  5.580 2.775 5.810 3.180 ;
        RECT  5.355 3.410 5.585 3.775 ;
        RECT  5.175 0.655 5.405 1.525 ;
        RECT  4.025 3.545 5.355 3.775 ;
        RECT  4.390 0.655 5.175 0.885 ;
        RECT  5.140 1.965 5.145 2.975 ;
        RECT  4.945 1.755 5.140 2.975 ;
        RECT  4.915 1.410 4.945 2.975 ;
        RECT  4.910 1.410 4.915 2.195 ;
        RECT  3.935 2.745 4.915 2.975 ;
        RECT  4.715 1.410 4.910 1.985 ;
        RECT  4.395 2.215 4.680 2.445 ;
        RECT  4.165 1.125 4.395 2.445 ;
        RECT  3.460 1.125 4.165 1.355 ;
        RECT  3.795 3.545 4.025 4.205 ;
        RECT  3.705 2.160 3.935 2.975 ;
        RECT  2.650 3.975 3.795 4.205 ;
        RECT  3.230 0.655 3.460 3.675 ;
        RECT  2.755 0.655 3.230 1.025 ;
        RECT  2.885 3.445 3.230 3.675 ;
        RECT  2.730 1.295 2.960 2.710 ;
        RECT  2.360 1.295 2.730 1.525 ;
        RECT  2.650 2.480 2.730 2.710 ;
        RECT  2.420 2.480 2.650 4.205 ;
        RECT  1.840 2.480 2.420 2.710 ;
        RECT  2.060 4.005 2.190 4.235 ;
        RECT  1.830 2.940 2.060 4.235 ;
        RECT  1.610 2.330 1.840 2.710 ;
        RECT  1.655 2.940 1.830 3.170 ;
        RECT  0.465 2.330 1.610 2.560 ;
        RECT  0.465 1.100 0.520 1.440 ;
        RECT  0.350 3.455 0.520 3.795 ;
        RECT  0.350 1.100 0.465 2.560 ;
        RECT  0.235 1.100 0.350 3.795 ;
        RECT  0.180 1.100 0.235 1.440 ;
        RECT  0.120 2.245 0.235 3.795 ;
    END
END DFFTRXL

MACRO DFFTRX4
    CLASS CORE ;
    FOREIGN DFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFTRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 1.250 1.940 1.590 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.550 1.260 15.700 2.660 ;
        RECT  15.465 1.260 15.550 3.020 ;
        RECT  15.320 0.805 15.465 3.020 ;
        RECT  15.125 0.805 15.320 1.615 ;
        RECT  15.235 2.790 15.320 3.020 ;
        RECT  15.005 2.790 15.235 3.625 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.740 0.805 13.970 1.620 ;
        RECT  13.720 2.890 13.850 3.230 ;
        RECT  13.720 1.260 13.740 1.620 ;
        RECT  13.510 1.260 13.720 3.230 ;
        RECT  13.490 1.260 13.510 3.120 ;
        RECT  13.340 1.260 13.490 2.660 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 1.820 2.500 2.300 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 1.820 1.355 2.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.185 -0.400 16.500 0.400 ;
        RECT  15.845 -0.400 16.185 0.950 ;
        RECT  14.745 -0.400 15.845 0.400 ;
        RECT  14.405 -0.400 14.745 1.420 ;
        RECT  13.305 -0.400 14.405 0.400 ;
        RECT  12.965 -0.400 13.305 0.950 ;
        RECT  12.000 -0.400 12.965 0.400 ;
        RECT  11.660 -0.400 12.000 0.575 ;
        RECT  9.265 -0.400 11.660 0.400 ;
        RECT  8.925 -0.400 9.265 1.215 ;
        RECT  6.660 -0.400 8.925 0.400 ;
        RECT  6.320 -0.400 6.660 1.190 ;
        RECT  4.440 -0.400 6.320 0.400 ;
        RECT  4.100 -0.400 4.440 1.270 ;
        RECT  1.240 -0.400 4.100 0.400 ;
        RECT  0.900 -0.400 1.240 0.950 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.050 4.640 16.500 5.440 ;
        RECT  15.710 3.445 16.050 5.440 ;
        RECT  14.570 4.640 15.710 5.440 ;
        RECT  14.230 4.040 14.570 5.440 ;
        RECT  13.130 4.640 14.230 5.440 ;
        RECT  12.790 4.070 13.130 5.440 ;
        RECT  11.830 4.640 12.790 5.440 ;
        RECT  11.490 4.465 11.830 5.440 ;
        RECT  9.215 4.640 11.490 5.440 ;
        RECT  8.985 3.570 9.215 5.440 ;
        RECT  5.900 4.640 8.985 5.440 ;
        RECT  5.845 4.465 5.900 5.440 ;
        RECT  5.615 4.410 5.845 5.440 ;
        RECT  5.560 4.465 5.615 5.440 ;
        RECT  4.310 4.640 5.560 5.440 ;
        RECT  3.970 4.465 4.310 5.440 ;
        RECT  1.285 4.640 3.970 5.440 ;
        RECT  0.945 3.760 1.285 5.440 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.860 2.030 15.090 2.375 ;
        RECT  14.775 2.145 14.860 2.375 ;
        RECT  14.545 2.145 14.775 3.690 ;
        RECT  12.755 3.460 14.545 3.690 ;
        RECT  12.755 1.310 12.765 1.650 ;
        RECT  12.525 1.310 12.755 3.690 ;
        RECT  12.425 1.310 12.525 1.650 ;
        RECT  12.250 3.150 12.525 3.490 ;
        RECT  12.065 2.015 12.295 2.370 ;
        RECT  11.445 3.205 12.250 3.435 ;
        RECT  11.990 2.015 12.065 2.245 ;
        RECT  11.760 1.405 11.990 2.245 ;
        RECT  10.545 1.405 11.760 1.635 ;
        RECT  11.215 3.205 11.445 3.610 ;
        RECT  10.955 1.885 11.170 2.115 ;
        RECT  10.725 1.885 10.955 4.335 ;
        RECT  9.885 4.105 10.725 4.335 ;
        RECT  10.495 1.250 10.545 1.635 ;
        RECT  10.265 1.250 10.495 3.270 ;
        RECT  10.205 1.250 10.265 1.675 ;
        RECT  8.295 2.605 10.265 2.835 ;
        RECT  8.225 1.445 10.205 1.675 ;
        RECT  9.655 3.075 9.885 4.335 ;
        RECT  8.755 3.075 9.655 3.305 ;
        RECT  8.525 3.075 8.755 3.735 ;
        RECT  7.355 3.505 8.525 3.735 ;
        RECT  8.065 2.605 8.295 3.115 ;
        RECT  7.995 1.145 8.225 1.675 ;
        RECT  7.935 2.885 8.065 3.115 ;
        RECT  7.640 1.145 7.995 1.375 ;
        RECT  7.705 2.885 7.935 3.240 ;
        RECT  7.355 2.390 7.835 2.620 ;
        RECT  7.125 2.390 7.355 3.735 ;
        RECT  5.600 3.505 7.125 3.735 ;
        RECT  6.665 1.420 6.895 3.100 ;
        RECT  6.020 1.420 6.665 1.650 ;
        RECT  5.830 2.870 6.665 3.100 ;
        RECT  6.325 2.190 6.435 2.530 ;
        RECT  6.095 1.880 6.325 2.530 ;
        RECT  5.160 1.880 6.095 2.110 ;
        RECT  5.790 1.160 6.020 1.650 ;
        RECT  5.625 1.160 5.790 1.390 ;
        RECT  5.600 2.340 5.765 2.570 ;
        RECT  5.395 0.630 5.625 1.390 ;
        RECT  5.370 2.340 5.600 3.735 ;
        RECT  5.190 0.630 5.395 0.860 ;
        RECT  4.990 3.505 5.370 3.735 ;
        RECT  5.140 1.350 5.160 2.110 ;
        RECT  4.910 1.350 5.140 2.935 ;
        RECT  4.760 3.505 4.990 4.165 ;
        RECT  4.820 1.350 4.910 1.690 ;
        RECT  3.770 2.705 4.910 2.935 ;
        RECT  2.675 3.935 4.760 4.165 ;
        RECT  4.450 1.980 4.680 2.320 ;
        RECT  3.420 1.980 4.450 2.210 ;
        RECT  3.190 0.745 3.420 3.515 ;
        RECT  2.740 0.745 3.190 0.975 ;
        RECT  3.135 3.285 3.190 3.515 ;
        RECT  2.905 3.285 3.135 3.690 ;
        RECT  2.730 1.360 2.960 2.785 ;
        RECT  2.655 1.360 2.730 1.590 ;
        RECT  2.675 2.535 2.730 2.785 ;
        RECT  2.445 2.535 2.675 4.165 ;
        RECT  2.425 1.240 2.655 1.590 ;
        RECT  0.520 2.535 2.445 2.765 ;
        RECT  1.985 3.015 2.215 4.100 ;
        RECT  1.500 3.015 1.985 3.245 ;
        RECT  0.415 0.745 0.520 1.555 ;
        RECT  0.415 2.535 0.520 4.045 ;
        RECT  0.185 0.745 0.415 4.045 ;
        RECT  0.180 0.745 0.185 1.555 ;
        RECT  0.180 2.765 0.185 4.045 ;
    END
END DFFTRX4

MACRO DFFTRX2
    CLASS CORE ;
    FOREIGN DFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFTRXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.845 1.765 2.435 ;
        RECT  1.260 2.205 1.460 2.435 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.625 2.635 13.680 4.025 ;
        RECT  13.625 1.285 13.645 1.515 ;
        RECT  13.565 1.285 13.625 4.025 ;
        RECT  13.395 0.810 13.565 4.025 ;
        RECT  13.225 0.810 13.395 1.620 ;
        RECT  13.340 2.745 13.395 4.025 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.185 2.405 12.325 2.635 ;
        RECT  12.125 0.960 12.185 3.080 ;
        RECT  11.955 0.905 12.125 3.080 ;
        RECT  11.785 0.905 11.955 1.245 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 0.725 2.425 0.955 ;
        RECT  2.035 0.725 2.265 1.590 ;
        RECT  1.715 1.360 2.035 1.590 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.990 1.285 1.105 1.515 ;
        RECT  0.760 1.285 0.990 2.335 ;
        RECT  0.645 1.980 0.760 2.335 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.845 -0.400 13.860 0.400 ;
        RECT  12.505 -0.400 12.845 1.420 ;
        RECT  10.700 -0.400 12.505 0.400 ;
        RECT  10.360 -0.400 10.700 1.100 ;
        RECT  8.640 -0.400 10.360 0.400 ;
        RECT  8.300 -0.400 8.640 1.225 ;
        RECT  5.985 -0.400 8.300 0.400 ;
        RECT  5.755 -0.400 5.985 0.945 ;
        RECT  4.125 -0.400 5.755 0.400 ;
        RECT  3.895 -0.400 4.125 0.870 ;
        RECT  1.080 -0.400 3.895 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.960 4.640 13.860 5.440 ;
        RECT  12.620 3.960 12.960 5.440 ;
        RECT  9.430 4.640 12.620 5.440 ;
        RECT  9.375 4.465 9.430 5.440 ;
        RECT  9.145 4.410 9.375 5.440 ;
        RECT  9.090 4.465 9.145 5.440 ;
        RECT  6.790 4.640 9.090 5.440 ;
        RECT  6.450 3.795 6.790 5.440 ;
        RECT  4.430 4.640 6.450 5.440 ;
        RECT  4.090 4.465 4.430 5.440 ;
        RECT  1.280 4.640 4.090 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.935 2.030 13.165 2.370 ;
        RECT  12.825 2.030 12.935 3.605 ;
        RECT  12.705 2.085 12.825 3.605 ;
        RECT  11.730 3.375 12.705 3.605 ;
        RECT  11.725 3.375 11.730 3.845 ;
        RECT  11.495 1.520 11.725 3.845 ;
        RECT  11.420 1.520 11.495 1.750 ;
        RECT  11.355 3.505 11.495 3.845 ;
        RECT  11.085 0.900 11.420 1.750 ;
        RECT  11.030 1.995 11.260 2.780 ;
        RECT  11.080 0.900 11.085 1.240 ;
        RECT  10.615 1.520 11.085 1.750 ;
        RECT  10.030 2.550 11.030 2.780 ;
        RECT  10.385 1.520 10.615 2.220 ;
        RECT  10.275 1.880 10.385 2.220 ;
        RECT  9.985 2.550 10.030 2.890 ;
        RECT  9.920 1.455 9.985 2.890 ;
        RECT  9.755 1.455 9.920 3.160 ;
        RECT  9.340 1.455 9.755 1.685 ;
        RECT  9.690 2.550 9.755 3.160 ;
        RECT  8.110 2.930 9.690 3.160 ;
        RECT  9.295 1.915 9.525 2.260 ;
        RECT  9.000 1.030 9.340 1.685 ;
        RECT  6.845 1.915 9.295 2.145 ;
        RECT  7.305 1.455 9.000 1.685 ;
        RECT  7.540 2.415 8.110 2.645 ;
        RECT  7.880 2.930 8.110 3.640 ;
        RECT  7.770 3.300 7.880 3.640 ;
        RECT  7.310 2.415 7.540 3.565 ;
        RECT  6.020 3.335 7.310 3.565 ;
        RECT  7.075 1.090 7.305 1.685 ;
        RECT  6.615 1.175 6.845 3.105 ;
        RECT  5.525 1.175 6.615 1.405 ;
        RECT  5.950 2.875 6.615 3.105 ;
        RECT  5.065 2.005 6.385 2.350 ;
        RECT  5.790 3.335 6.020 4.055 ;
        RECT  3.670 3.825 5.790 4.055 ;
        RECT  5.295 0.885 5.525 1.405 ;
        RECT  5.185 0.885 5.295 1.115 ;
        RECT  4.955 0.630 5.185 1.115 ;
        RECT  4.835 1.590 5.065 3.365 ;
        RECT  4.370 0.630 4.955 0.860 ;
        RECT  4.640 1.590 4.835 1.820 ;
        RECT  4.020 3.135 4.835 3.365 ;
        RECT  4.375 2.110 4.605 2.525 ;
        RECT  3.190 2.295 4.375 2.525 ;
        RECT  3.790 2.780 4.020 3.365 ;
        RECT  3.680 2.780 3.790 3.120 ;
        RECT  3.440 3.825 3.670 4.155 ;
        RECT  2.595 3.925 3.440 4.155 ;
        RECT  3.185 1.010 3.190 2.525 ;
        RECT  3.055 1.010 3.185 2.965 ;
        RECT  2.960 1.010 3.055 3.650 ;
        RECT  2.955 0.895 2.960 3.650 ;
        RECT  2.730 0.895 2.955 1.240 ;
        RECT  2.825 2.735 2.955 3.650 ;
        RECT  2.595 1.820 2.725 2.050 ;
        RECT  2.365 1.820 2.595 4.155 ;
        RECT  0.520 2.665 2.365 2.895 ;
        RECT  1.905 3.125 2.135 4.210 ;
        RECT  1.540 3.125 1.905 3.355 ;
        RECT  0.415 1.310 0.520 1.650 ;
        RECT  0.415 2.665 0.520 3.530 ;
        RECT  0.185 1.310 0.415 3.530 ;
        RECT  0.180 1.310 0.185 1.650 ;
        RECT  0.180 3.190 0.185 3.530 ;
    END
END DFFTRX2

MACRO DFFTRX1
    CLASS CORE ;
    FOREIGN DFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFTRXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 1.710 1.840 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.865 1.845 11.005 2.075 ;
        RECT  10.810 1.200 10.865 2.075 ;
        RECT  10.635 1.200 10.810 3.230 ;
        RECT  10.580 1.845 10.635 3.230 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 0.805 10.345 3.800 ;
        RECT  9.365 0.805 10.115 1.035 ;
        RECT  9.445 3.570 10.115 3.800 ;
        RECT  9.105 3.570 9.445 3.910 ;
        RECT  9.135 0.660 9.365 1.035 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.070 1.895 2.500 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 2.790 1.230 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.160 -0.400 11.220 0.400 ;
        RECT  9.820 -0.400 10.160 0.575 ;
        RECT  8.700 -0.400 9.820 0.400 ;
        RECT  8.360 -0.400 8.700 0.950 ;
        RECT  5.965 -0.400 8.360 0.400 ;
        RECT  5.735 -0.400 5.965 0.900 ;
        RECT  4.105 -0.400 5.735 0.400 ;
        RECT  3.875 -0.400 4.105 0.870 ;
        RECT  0.600 -0.400 3.875 0.400 ;
        RECT  0.260 -0.400 0.600 0.575 ;
        RECT  0.000 -0.400 0.260 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.145 4.640 11.220 5.440 ;
        RECT  10.090 4.465 10.145 5.440 ;
        RECT  9.860 4.410 10.090 5.440 ;
        RECT  9.805 4.465 9.860 5.440 ;
        RECT  8.725 4.640 9.805 5.440 ;
        RECT  8.385 3.960 8.725 5.440 ;
        RECT  6.365 4.640 8.385 5.440 ;
        RECT  6.025 3.540 6.365 5.440 ;
        RECT  4.620 4.640 6.025 5.440 ;
        RECT  4.565 4.465 4.620 5.440 ;
        RECT  4.335 4.410 4.565 5.440 ;
        RECT  4.280 4.465 4.335 5.440 ;
        RECT  1.315 4.640 4.280 5.440 ;
        RECT  0.905 4.465 1.315 5.440 ;
        RECT  0.000 4.640 0.905 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.545 1.490 9.885 3.130 ;
        RECT  9.120 1.490 9.545 1.830 ;
        RECT  9.105 2.790 9.545 3.130 ;
        RECT  8.275 1.520 9.120 1.750 ;
        RECT  8.870 2.140 9.090 2.480 ;
        RECT  8.750 2.140 8.870 2.725 ;
        RECT  8.640 2.250 8.750 2.725 ;
        RECT  7.670 2.495 8.640 2.725 ;
        RECT  8.045 1.520 8.275 2.220 ;
        RECT  7.670 3.600 7.725 3.940 ;
        RECT  7.440 1.215 7.670 3.940 ;
        RECT  7.285 1.215 7.440 1.445 ;
        RECT  7.385 3.600 7.440 3.940 ;
        RECT  7.055 1.090 7.285 1.445 ;
        RECT  6.825 1.885 7.100 2.115 ;
        RECT  6.595 1.295 6.825 3.005 ;
        RECT  5.370 1.295 6.595 1.525 ;
        RECT  5.810 2.775 6.595 3.005 ;
        RECT  5.145 1.965 6.365 2.345 ;
        RECT  5.580 2.775 5.810 3.180 ;
        RECT  5.355 3.410 5.585 3.775 ;
        RECT  5.135 0.655 5.370 1.525 ;
        RECT  4.025 3.545 5.355 3.775 ;
        RECT  5.140 1.965 5.145 2.975 ;
        RECT  4.915 1.755 5.140 2.975 ;
        RECT  4.350 0.655 5.135 0.885 ;
        RECT  4.910 1.755 4.915 2.195 ;
        RECT  3.895 2.745 4.915 2.975 ;
        RECT  4.905 1.755 4.910 1.985 ;
        RECT  4.675 1.410 4.905 1.985 ;
        RECT  4.355 2.215 4.680 2.445 ;
        RECT  4.125 1.125 4.355 2.445 ;
        RECT  3.385 1.125 4.125 1.355 ;
        RECT  3.795 3.545 4.025 4.205 ;
        RECT  3.665 2.160 3.895 2.975 ;
        RECT  2.650 3.975 3.795 4.205 ;
        RECT  3.155 0.655 3.385 3.675 ;
        RECT  2.715 0.655 3.155 1.025 ;
        RECT  2.885 3.445 3.155 3.675 ;
        RECT  2.405 1.375 2.660 1.605 ;
        RECT  2.420 2.890 2.650 4.205 ;
        RECT  1.840 2.890 2.420 3.120 ;
        RECT  2.175 0.875 2.405 1.605 ;
        RECT  2.060 4.150 2.190 4.380 ;
        RECT  0.520 0.875 2.175 1.105 ;
        RECT  1.830 3.350 2.060 4.380 ;
        RECT  1.610 2.330 1.840 3.120 ;
        RECT  1.655 3.350 1.830 3.580 ;
        RECT  0.465 2.330 1.610 2.560 ;
        RECT  0.465 0.875 0.520 1.500 ;
        RECT  0.350 3.450 0.520 3.680 ;
        RECT  0.350 0.875 0.465 2.560 ;
        RECT  0.290 0.875 0.350 3.680 ;
        RECT  0.235 1.160 0.290 3.680 ;
        RECT  0.180 1.160 0.235 1.500 ;
        RECT  0.120 2.245 0.235 3.680 ;
    END
END DFFTRX1

MACRO DFFSRHQXL
    CLASS CORE ;
    FOREIGN DFFSRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.785 2.885 15.125 3.225 ;
        RECT  14.075 2.940 14.785 3.170 ;
        RECT  13.930 2.940 14.075 3.220 ;
        RECT  13.930 2.250 13.985 2.590 ;
        RECT  13.700 2.250 13.930 4.045 ;
        RECT  13.645 2.250 13.700 2.590 ;
        RECT  10.470 3.815 13.700 4.045 ;
        RECT  10.430 2.765 10.470 4.045 ;
        RECT  10.420 2.710 10.430 4.045 ;
        RECT  10.345 2.660 10.420 4.045 ;
        RECT  10.240 2.405 10.345 4.045 ;
        RECT  10.090 2.405 10.240 3.240 ;
        RECT  9.510 3.010 10.090 3.240 ;
        RECT  9.280 3.010 9.510 4.405 ;
        RECT  6.820 4.175 9.280 4.405 ;
        RECT  6.590 3.445 6.820 4.405 ;
        RECT  5.895 3.445 6.590 3.675 ;
        RECT  5.665 3.445 5.895 4.410 ;
        RECT  3.990 4.180 5.665 4.410 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.850 2.405 12.985 2.635 ;
        RECT  12.230 2.315 12.850 2.855 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.600 1.845 15.625 2.075 ;
        RECT  15.370 1.330 15.600 3.945 ;
        RECT  14.560 1.330 15.370 1.560 ;
        RECT  14.890 3.715 15.370 3.945 ;
        RECT  14.550 3.660 14.890 4.000 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.850 2.060 1.400 2.765 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 3.810 0.625 4.150 ;
        RECT  0.150 3.810 0.620 4.390 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.450 -0.400 15.840 0.400 ;
        RECT  13.110 -0.400 13.450 1.555 ;
        RECT  9.790 -0.400 13.110 0.400 ;
        RECT  9.450 -0.400 9.790 0.575 ;
        RECT  7.110 -0.400 9.450 0.400 ;
        RECT  6.770 -0.400 7.110 1.075 ;
        RECT  3.665 -0.400 6.770 0.400 ;
        RECT  3.325 -0.400 3.665 0.900 ;
        RECT  1.205 -0.400 3.325 0.400 ;
        RECT  0.865 -0.400 1.205 0.575 ;
        RECT  0.000 -0.400 0.865 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.660 4.640 15.840 5.440 ;
        RECT  15.320 4.465 15.660 5.440 ;
        RECT  13.550 4.640 15.320 5.440 ;
        RECT  13.210 4.465 13.550 5.440 ;
        RECT  12.345 4.640 13.210 5.440 ;
        RECT  12.005 4.465 12.345 5.440 ;
        RECT  10.010 4.640 12.005 5.440 ;
        RECT  9.780 3.640 10.010 5.440 ;
        RECT  6.355 4.640 9.780 5.440 ;
        RECT  6.125 3.915 6.355 5.440 ;
        RECT  3.660 4.640 6.125 5.440 ;
        RECT  3.320 4.465 3.660 5.440 ;
        RECT  1.195 4.640 3.320 5.440 ;
        RECT  0.855 4.465 1.195 5.440 ;
        RECT  0.000 4.640 0.855 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.510 0.870 15.660 1.100 ;
        RECT  15.280 0.795 15.510 1.100 ;
        RECT  14.170 0.795 15.280 1.025 ;
        RECT  14.980 1.970 15.090 2.310 ;
        RECT  14.750 1.790 14.980 2.310 ;
        RECT  12.690 1.790 14.750 2.020 ;
        RECT  13.940 0.795 14.170 1.555 ;
        RECT  13.830 1.215 13.940 1.555 ;
        RECT  13.405 2.975 13.460 3.205 ;
        RECT  13.120 2.975 13.405 3.525 ;
        RECT  11.885 3.295 13.120 3.525 ;
        RECT  12.350 1.420 12.690 2.020 ;
        RECT  11.885 1.790 12.350 2.020 ;
        RECT  12.000 0.775 12.190 1.005 ;
        RECT  11.770 0.775 12.000 1.505 ;
        RECT  11.655 1.790 11.885 3.525 ;
        RECT  10.250 1.275 11.770 1.505 ;
        RECT  11.335 1.740 11.390 1.970 ;
        RECT  10.930 1.735 11.335 1.980 ;
        RECT  10.775 0.660 11.005 1.035 ;
        RECT  10.700 1.735 10.930 3.580 ;
        RECT  9.910 0.805 10.775 1.035 ;
        RECT  9.530 1.750 10.700 2.015 ;
        RECT  9.680 0.805 9.910 1.270 ;
        RECT  9.045 1.040 9.680 1.270 ;
        RECT  9.295 1.750 9.530 2.120 ;
        RECT  8.815 1.040 9.045 3.170 ;
        RECT  8.645 3.605 8.985 3.945 ;
        RECT  8.290 1.040 8.815 1.270 ;
        RECT  8.560 2.940 8.815 3.170 ;
        RECT  7.280 3.715 8.645 3.945 ;
        RECT  8.350 1.500 8.580 2.710 ;
        RECT  8.220 2.940 8.560 3.280 ;
        RECT  7.910 1.500 8.350 1.730 ;
        RECT  7.740 2.480 8.350 2.710 ;
        RECT  7.280 1.960 8.115 2.190 ;
        RECT  7.680 1.070 7.910 1.730 ;
        RECT  7.510 2.480 7.740 3.480 ;
        RECT  7.570 1.070 7.680 1.410 ;
        RECT  7.050 1.310 7.280 3.945 ;
        RECT  6.310 1.310 7.050 1.540 ;
        RECT  6.075 2.975 7.050 3.205 ;
        RECT  6.465 2.200 6.780 2.540 ;
        RECT  6.440 1.775 6.465 2.540 ;
        RECT  6.235 1.775 6.440 2.485 ;
        RECT  6.150 1.200 6.310 1.540 ;
        RECT  5.005 1.775 6.235 2.005 ;
        RECT  5.970 0.630 6.150 1.540 ;
        RECT  5.920 0.630 5.970 1.485 ;
        RECT  5.615 2.240 5.955 2.580 ;
        RECT  5.810 0.630 5.920 0.970 ;
        RECT  5.430 2.350 5.615 2.580 ;
        RECT  5.200 2.350 5.430 3.845 ;
        RECT  2.840 3.615 5.200 3.845 ;
        RECT  4.970 1.300 5.005 2.005 ;
        RECT  4.740 1.300 4.970 3.325 ;
        RECT  4.665 1.300 4.740 1.640 ;
        RECT  3.400 3.095 4.740 3.325 ;
        RECT  4.280 2.005 4.510 2.380 ;
        RECT  2.625 2.005 4.280 2.235 ;
        RECT  3.170 2.525 3.400 3.325 ;
        RECT  3.050 2.525 3.170 2.755 ;
        RECT  2.610 3.615 2.840 4.345 ;
        RECT  2.440 1.195 2.625 2.735 ;
        RECT  1.885 4.115 2.610 4.345 ;
        RECT  2.395 1.140 2.440 2.735 ;
        RECT  2.100 1.140 2.395 1.480 ;
        RECT  2.345 2.505 2.395 2.735 ;
        RECT  2.115 2.505 2.345 3.825 ;
        RECT  1.885 1.825 2.150 2.055 ;
        RECT  1.655 1.825 1.885 4.345 ;
        RECT  0.520 3.220 1.655 3.450 ;
        RECT  0.465 1.210 0.520 1.550 ;
        RECT  0.465 3.165 0.520 3.505 ;
        RECT  0.235 1.210 0.465 3.505 ;
        RECT  0.180 1.210 0.235 1.550 ;
        RECT  0.180 3.165 0.235 3.505 ;
    END
END DFFSRHQXL

MACRO DFFSRHQX4
    CLASS CORE ;
    FOREIGN DFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRHQXL ;
    SIZE 30.360 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.425 2.495 28.190 2.725 ;
        RECT  22.975 2.085 23.425 2.725 ;
        RECT  22.835 2.495 22.975 2.725 ;
        RECT  22.605 2.495 22.835 4.005 ;
        RECT  19.075 3.775 22.605 4.005 ;
        RECT  18.845 3.420 19.075 4.005 ;
        RECT  17.710 3.420 18.845 3.650 ;
        RECT  17.710 2.315 17.760 2.655 ;
        RECT  17.475 2.315 17.710 3.650 ;
        RECT  17.420 2.315 17.475 2.685 ;
        RECT  17.300 3.195 17.475 3.650 ;
        RECT  17.375 2.405 17.420 2.685 ;
        RECT  17.135 3.420 17.300 3.650 ;
        RECT  16.905 3.420 17.135 4.155 ;
        RECT  9.180 3.925 16.905 4.155 ;
        RECT  8.950 3.580 9.180 4.155 ;
        RECT  7.795 3.580 8.950 3.810 ;
        RECT  7.565 3.580 7.795 4.015 ;
        RECT  5.330 3.785 7.565 4.015 ;
        RECT  5.100 3.785 5.330 4.205 ;
        RECT  4.790 3.975 5.100 4.205 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.245 2.315 20.935 2.545 ;
        RECT  20.015 2.315 20.245 2.635 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  30.145 2.380 30.220 3.780 ;
        RECT  30.070 2.075 30.145 3.780 ;
        RECT  29.840 1.370 30.070 3.780 ;
        RECT  29.460 1.370 29.840 1.600 ;
        RECT  29.150 2.960 29.840 3.600 ;
        RECT  28.825 1.260 29.460 1.600 ;
        RECT  28.050 2.960 29.150 3.295 ;
        RECT  28.020 1.315 28.825 1.600 ;
        RECT  27.765 2.960 28.050 3.835 ;
        RECT  27.505 1.260 28.020 1.600 ;
        RECT  27.710 3.025 27.765 3.835 ;
        RECT  26.260 3.065 27.710 3.295 ;
        RECT  26.615 1.370 27.505 1.600 ;
        RECT  26.240 1.260 26.615 1.600 ;
        RECT  26.050 3.065 26.260 3.530 ;
        RECT  25.710 2.975 26.050 3.795 ;
        RECT  23.620 3.110 25.710 3.340 ;
        RECT  23.410 3.110 23.620 3.530 ;
        RECT  23.070 3.060 23.410 3.880 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 2.210 1.905 2.550 ;
        RECT  1.460 2.210 1.845 2.910 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.755 2.090 0.760 2.375 ;
        RECT  0.375 1.880 0.755 2.660 ;
        RECT  0.215 2.100 0.375 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.160 -0.400 30.360 0.400 ;
        RECT  24.820 -0.400 25.160 0.895 ;
        RECT  23.675 -0.400 24.820 0.400 ;
        RECT  23.335 -0.400 23.675 0.895 ;
        RECT  22.100 -0.400 23.335 0.400 ;
        RECT  21.760 -0.400 22.100 1.335 ;
        RECT  20.555 -0.400 21.760 0.400 ;
        RECT  20.555 1.200 20.580 1.540 ;
        RECT  20.325 -0.400 20.555 1.540 ;
        RECT  17.475 -0.400 20.325 0.400 ;
        RECT  20.240 1.200 20.325 1.540 ;
        RECT  17.135 -0.400 17.475 0.575 ;
        RECT  12.290 -0.400 17.135 0.400 ;
        RECT  11.950 -0.400 12.290 0.815 ;
        RECT  10.755 -0.400 11.950 0.400 ;
        RECT  10.415 -0.400 10.755 0.815 ;
        RECT  9.830 -0.400 10.415 0.400 ;
        RECT  9.490 -0.400 9.830 1.090 ;
        RECT  5.565 -0.400 9.490 0.400 ;
        RECT  4.285 -0.400 5.565 0.870 ;
        RECT  1.500 -0.400 4.285 0.400 ;
        RECT  1.160 -0.400 1.500 0.575 ;
        RECT  0.000 -0.400 1.160 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  28.770 4.640 30.360 5.440 ;
        RECT  28.430 3.530 28.770 5.440 ;
        RECT  27.330 4.640 28.430 5.440 ;
        RECT  26.990 3.530 27.330 5.440 ;
        RECT  24.730 4.640 26.990 5.440 ;
        RECT  24.390 3.740 24.730 5.440 ;
        RECT  21.770 4.640 24.390 5.440 ;
        RECT  21.430 4.465 21.770 5.440 ;
        RECT  20.185 4.640 21.430 5.440 ;
        RECT  19.845 4.465 20.185 5.440 ;
        RECT  17.705 4.640 19.845 5.440 ;
        RECT  17.365 3.880 17.705 5.440 ;
        RECT  8.365 4.640 17.365 5.440 ;
        RECT  8.025 4.090 8.365 5.440 ;
        RECT  6.035 4.640 8.025 5.440 ;
        RECT  5.695 4.465 6.035 5.440 ;
        RECT  4.540 4.640 5.695 5.440 ;
        RECT  4.310 3.755 4.540 5.440 ;
        RECT  1.825 4.640 4.310 5.440 ;
        RECT  1.485 3.645 1.825 5.440 ;
        RECT  0.000 4.640 1.485 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  29.840 0.710 30.180 1.050 ;
        RECT  28.740 0.765 29.840 0.995 ;
        RECT  28.950 1.960 29.290 2.300 ;
        RECT  23.980 2.015 28.950 2.245 ;
        RECT  28.400 0.690 28.740 1.030 ;
        RECT  27.300 0.745 28.400 0.975 ;
        RECT  26.960 0.690 27.300 1.030 ;
        RECT  25.860 0.745 26.960 0.975 ;
        RECT  25.630 0.745 25.860 1.355 ;
        RECT  25.520 1.015 25.630 1.355 ;
        RECT  24.435 1.125 25.520 1.355 ;
        RECT  24.095 0.945 24.435 1.355 ;
        RECT  22.955 1.125 24.095 1.355 ;
        RECT  23.750 1.585 23.980 2.245 ;
        RECT  22.370 1.585 23.750 1.815 ;
        RECT  22.615 1.015 22.955 1.355 ;
        RECT  22.140 1.585 22.370 2.590 ;
        RECT  21.405 2.360 22.140 2.590 ;
        RECT  21.400 1.375 21.405 2.590 ;
        RECT  21.300 1.375 21.400 3.420 ;
        RECT  21.170 1.320 21.300 3.420 ;
        RECT  20.960 1.320 21.170 1.660 ;
        RECT  20.970 3.190 21.170 3.420 ;
        RECT  20.630 3.190 20.970 3.530 ;
        RECT  19.590 3.245 20.630 3.475 ;
        RECT  19.595 0.750 19.825 1.425 ;
        RECT  19.590 2.180 19.645 2.520 ;
        RECT  18.495 0.750 19.595 0.980 ;
        RECT  19.360 2.180 19.590 3.475 ;
        RECT  19.305 2.180 19.360 2.520 ;
        RECT  18.845 1.215 19.075 2.655 ;
        RECT  18.735 1.215 18.845 1.620 ;
        RECT  18.250 2.425 18.845 2.655 ;
        RECT  17.005 1.390 18.735 1.620 ;
        RECT  16.400 1.850 18.585 2.080 ;
        RECT  18.265 0.750 18.495 1.155 ;
        RECT  17.935 0.925 18.265 1.155 ;
        RECT  18.020 2.425 18.250 3.190 ;
        RECT  16.775 1.215 17.005 1.620 ;
        RECT  16.445 2.355 16.675 3.620 ;
        RECT  15.855 2.355 16.445 2.585 ;
        RECT  16.175 3.390 16.445 3.620 ;
        RECT  16.170 0.770 16.400 2.080 ;
        RECT  15.190 2.905 16.215 3.135 ;
        RECT  15.805 3.390 16.175 3.675 ;
        RECT  16.100 0.770 16.170 1.000 ;
        RECT  15.760 0.660 16.100 1.000 ;
        RECT  15.855 1.330 15.910 1.670 ;
        RECT  15.625 1.330 15.855 2.585 ;
        RECT  9.690 3.445 15.805 3.675 ;
        RECT  15.250 0.715 15.760 0.945 ;
        RECT  15.570 1.330 15.625 1.670 ;
        RECT  15.250 1.245 15.305 1.585 ;
        RECT  15.190 0.715 15.250 1.585 ;
        RECT  14.960 0.715 15.190 3.135 ;
        RECT  13.855 0.715 14.960 0.945 ;
        RECT  13.290 2.905 14.960 3.135 ;
        RECT  14.525 1.270 14.580 1.610 ;
        RECT  14.295 1.270 14.525 2.295 ;
        RECT  14.240 1.270 14.295 1.610 ;
        RECT  13.050 2.065 14.295 2.295 ;
        RECT  13.625 0.715 13.855 1.795 ;
        RECT  13.515 0.985 13.625 1.795 ;
        RECT  12.945 0.985 13.050 2.295 ;
        RECT  12.715 0.985 12.945 3.135 ;
        RECT  12.710 0.985 12.715 1.800 ;
        RECT  9.920 2.905 12.715 3.135 ;
        RECT  11.515 1.570 12.710 1.800 ;
        RECT  11.230 0.985 11.515 1.800 ;
        RECT  11.175 0.985 11.230 1.795 ;
        RECT  10.485 1.385 10.715 2.650 ;
        RECT  8.860 1.385 10.485 1.615 ;
        RECT  9.690 2.420 10.485 2.650 ;
        RECT  9.225 1.925 10.215 2.155 ;
        RECT  9.460 2.420 9.690 3.675 ;
        RECT  8.645 3.120 9.460 3.350 ;
        RECT  8.995 1.925 9.225 2.800 ;
        RECT  7.335 2.570 8.995 2.800 ;
        RECT  8.630 0.630 8.860 1.615 ;
        RECT  7.795 2.055 8.765 2.285 ;
        RECT  8.515 0.630 8.630 0.860 ;
        RECT  8.030 0.635 8.260 1.275 ;
        RECT  6.415 0.635 8.030 0.865 ;
        RECT  7.565 1.100 7.795 2.285 ;
        RECT  6.875 1.100 7.565 1.330 ;
        RECT  7.105 1.560 7.335 3.525 ;
        RECT  4.205 3.295 7.105 3.525 ;
        RECT  6.645 1.100 6.875 3.005 ;
        RECT  4.765 2.775 6.645 3.005 ;
        RECT  6.185 0.635 6.415 1.600 ;
        RECT  6.300 2.140 6.410 2.480 ;
        RECT  6.070 1.890 6.300 2.480 ;
        RECT  5.070 1.315 6.185 1.545 ;
        RECT  3.175 1.890 6.070 2.120 ;
        RECT  4.730 1.315 5.070 1.655 ;
        RECT  4.535 2.400 4.765 3.005 ;
        RECT  3.635 2.400 4.535 2.630 ;
        RECT  3.975 2.860 4.205 3.525 ;
        RECT  3.865 2.860 3.975 3.200 ;
        RECT  3.405 2.400 3.635 4.230 ;
        RECT  2.585 4.000 3.405 4.230 ;
        RECT  2.945 1.055 3.175 3.695 ;
        RECT  2.905 1.055 2.945 1.285 ;
        RECT  2.565 0.945 2.905 1.285 ;
        RECT  2.355 3.155 2.585 4.230 ;
        RECT  2.405 1.760 2.580 1.990 ;
        RECT  2.175 1.750 2.405 1.990 ;
        RECT  1.225 3.155 2.355 3.385 ;
        RECT  1.225 1.750 2.175 1.980 ;
        RECT  0.995 1.280 1.225 3.385 ;
        RECT  0.670 1.280 0.995 1.510 ;
        RECT  0.990 2.945 0.995 3.385 ;
        RECT  0.650 2.945 0.990 4.225 ;
        RECT  0.330 0.695 0.670 1.515 ;
    END
END DFFSRHQX4

MACRO DFFSRHQX2
    CLASS CORE ;
    FOREIGN DFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRHQXL ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 2.495 19.935 2.725 ;
        RECT  17.125 2.375 17.605 2.725 ;
        RECT  16.895 2.375 17.125 4.005 ;
        RECT  16.870 2.375 16.895 2.605 ;
        RECT  16.715 3.755 16.895 4.005 ;
        RECT  13.570 3.775 16.715 4.005 ;
        RECT  13.570 2.610 13.730 2.840 ;
        RECT  13.340 2.610 13.570 4.005 ;
        RECT  12.515 2.610 13.340 2.840 ;
        RECT  12.285 2.610 12.515 4.315 ;
        RECT  12.095 3.955 12.285 4.315 ;
        RECT  7.620 3.955 12.095 4.185 ;
        RECT  7.390 3.500 7.620 4.185 ;
        RECT  6.700 3.500 7.390 3.730 ;
        RECT  6.470 3.500 6.700 4.290 ;
        RECT  4.685 4.060 6.470 4.290 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.630 1.725 15.670 2.695 ;
        RECT  15.350 1.685 15.630 2.695 ;
        RECT  15.290 1.685 15.350 2.025 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.565 1.370 21.570 3.195 ;
        RECT  21.340 1.370 21.565 3.205 ;
        RECT  21.275 1.370 21.340 1.600 ;
        RECT  21.335 2.965 21.340 3.205 ;
        RECT  20.200 2.975 21.335 3.205 ;
        RECT  20.905 1.260 21.275 1.600 ;
        RECT  20.015 1.370 20.905 1.600 ;
        RECT  19.860 2.975 20.200 4.170 ;
        RECT  19.405 1.260 20.015 1.600 ;
        RECT  18.130 2.975 19.860 3.205 ;
        RECT  17.845 2.975 18.130 4.010 ;
        RECT  17.790 3.190 17.845 4.010 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 1.810 1.880 2.725 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 2.065 0.605 2.780 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.265 -0.400 22.440 0.400 ;
        RECT  17.925 -0.400 18.265 1.220 ;
        RECT  16.200 -0.400 17.925 0.400 ;
        RECT  15.860 -0.400 16.200 1.325 ;
        RECT  13.175 -0.400 15.860 0.400 ;
        RECT  12.835 -0.400 13.175 0.575 ;
        RECT  9.200 -0.400 12.835 0.400 ;
        RECT  8.860 -0.400 9.200 0.815 ;
        RECT  7.730 -0.400 8.860 0.400 ;
        RECT  7.390 -0.400 7.730 0.820 ;
        RECT  4.345 -0.400 7.390 0.400 ;
        RECT  4.005 -0.400 4.345 1.595 ;
        RECT  1.640 -0.400 4.005 0.400 ;
        RECT  1.300 -0.400 1.640 1.430 ;
        RECT  0.000 -0.400 1.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.920 4.640 22.440 5.440 ;
        RECT  20.580 3.615 20.920 5.440 ;
        RECT  19.480 4.640 20.580 5.440 ;
        RECT  19.140 3.595 19.480 5.440 ;
        RECT  16.760 4.640 19.140 5.440 ;
        RECT  16.420 4.465 16.760 5.440 ;
        RECT  15.350 4.640 16.420 5.440 ;
        RECT  15.010 4.465 15.350 5.440 ;
        RECT  13.105 4.640 15.010 5.440 ;
        RECT  12.875 3.600 13.105 5.440 ;
        RECT  7.160 4.640 12.875 5.440 ;
        RECT  6.930 3.960 7.160 5.440 ;
        RECT  4.425 4.640 6.930 5.440 ;
        RECT  4.195 3.960 4.425 5.440 ;
        RECT  1.610 4.640 4.195 5.440 ;
        RECT  1.270 3.650 1.610 5.440 ;
        RECT  0.000 4.640 1.270 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.035 1.125 22.145 1.465 ;
        RECT  21.805 0.800 22.035 1.465 ;
        RECT  20.510 0.800 21.805 1.030 ;
        RECT  20.875 1.915 21.105 2.350 ;
        RECT  16.925 1.915 20.875 2.145 ;
        RECT  20.170 0.690 20.510 1.030 ;
        RECT  19.025 0.800 20.170 1.030 ;
        RECT  18.970 0.800 19.025 1.490 ;
        RECT  18.795 0.800 18.970 1.685 ;
        RECT  18.685 1.150 18.795 1.685 ;
        RECT  17.465 1.455 18.685 1.685 ;
        RECT  17.235 0.750 17.465 1.685 ;
        RECT  17.125 0.750 17.235 1.090 ;
        RECT  16.585 1.455 16.925 2.145 ;
        RECT  16.520 1.915 16.585 2.145 ;
        RECT  16.410 1.915 16.520 2.755 ;
        RECT  16.290 1.915 16.410 3.255 ;
        RECT  16.180 2.415 16.290 3.255 ;
        RECT  16.110 3.025 16.180 3.255 ;
        RECT  15.770 3.025 16.110 3.365 ;
        RECT  15.105 3.025 15.770 3.255 ;
        RECT  15.250 1.150 15.500 1.380 ;
        RECT  15.020 0.825 15.250 1.380 ;
        RECT  14.875 2.420 15.105 3.255 ;
        RECT  13.540 0.825 15.020 1.055 ;
        RECT  14.695 2.420 14.875 2.650 ;
        RECT  14.625 1.345 14.680 1.575 ;
        RECT  14.435 1.285 14.625 1.575 ;
        RECT  14.205 1.285 14.435 3.300 ;
        RECT  12.835 1.285 14.205 1.515 ;
        RECT  14.030 3.070 14.205 3.300 ;
        RECT  13.800 3.070 14.030 3.460 ;
        RECT  13.745 1.850 13.975 2.325 ;
        RECT  11.750 2.095 13.745 2.325 ;
        RECT  12.605 1.285 12.835 1.860 ;
        RECT  12.495 1.520 12.605 1.860 ;
        RECT  11.380 3.330 12.050 3.560 ;
        RECT  11.675 2.795 11.995 3.025 ;
        RECT  11.750 0.690 11.805 0.920 ;
        RECT  11.675 0.690 11.750 2.325 ;
        RECT  11.445 0.690 11.675 3.025 ;
        RECT  10.645 0.795 11.445 1.025 ;
        RECT  10.710 2.795 11.445 3.025 ;
        RECT  11.150 3.330 11.380 3.645 ;
        RECT  10.980 1.460 11.210 2.045 ;
        RECT  8.080 3.415 11.150 3.645 ;
        RECT  9.860 1.815 10.980 2.045 ;
        RECT  10.370 2.740 10.710 3.080 ;
        RECT  10.415 0.795 10.645 1.585 ;
        RECT  10.195 1.355 10.415 1.585 ;
        RECT  9.790 0.750 10.085 0.980 ;
        RECT  9.600 2.740 9.940 3.080 ;
        RECT  9.470 1.515 9.860 2.045 ;
        RECT  9.560 0.750 9.790 1.280 ;
        RECT  8.540 2.795 9.600 3.025 ;
        RECT  7.865 1.050 9.560 1.280 ;
        RECT  8.540 1.815 9.470 2.045 ;
        RECT  8.310 1.515 8.540 3.080 ;
        RECT  8.095 1.515 8.310 1.745 ;
        RECT  7.865 3.015 8.080 3.645 ;
        RECT  7.850 1.050 7.865 3.645 ;
        RECT  7.635 1.050 7.850 3.245 ;
        RECT  6.930 1.255 7.635 1.485 ;
        RECT  6.940 3.015 7.635 3.245 ;
        RECT  7.175 1.770 7.405 2.520 ;
        RECT  5.775 1.770 7.175 2.000 ;
        RECT  6.820 1.200 6.930 1.540 ;
        RECT  6.590 0.655 6.820 1.540 ;
        RECT  6.235 2.235 6.755 2.465 ;
        RECT  6.420 0.655 6.590 0.885 ;
        RECT  6.005 2.235 6.235 3.675 ;
        RECT  3.470 3.445 6.005 3.675 ;
        RECT  5.665 1.445 5.775 3.215 ;
        RECT  5.545 1.390 5.665 3.215 ;
        RECT  5.325 1.390 5.545 1.730 ;
        RECT  4.415 2.985 5.545 3.215 ;
        RECT  3.015 2.115 5.310 2.345 ;
        RECT  4.185 2.595 4.415 3.215 ;
        RECT  3.860 2.595 4.185 2.825 ;
        RECT  3.240 3.030 3.470 4.410 ;
        RECT  2.540 4.170 3.240 4.410 ;
        RECT  3.005 1.225 3.015 2.345 ;
        RECT  2.980 1.225 3.005 3.910 ;
        RECT  2.775 1.170 2.980 3.910 ;
        RECT  2.640 1.170 2.775 1.510 ;
        RECT  2.500 3.045 2.540 4.410 ;
        RECT  2.270 1.930 2.500 4.410 ;
        RECT  1.070 3.045 2.270 3.275 ;
        RECT  0.870 1.200 1.070 3.275 ;
        RECT  0.840 1.145 0.870 3.275 ;
        RECT  0.530 1.145 0.840 1.485 ;
        RECT  0.730 3.045 0.840 3.275 ;
        RECT  0.445 3.045 0.730 4.195 ;
        RECT  0.390 3.375 0.445 4.195 ;
    END
END DFFSRHQX2

MACRO DFFSRHQX1
    CLASS CORE ;
    FOREIGN DFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRHQXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.910 2.610 15.140 2.950 ;
        RECT  13.930 2.665 14.910 2.895 ;
        RECT  13.700 2.250 13.930 4.235 ;
        RECT  10.470 4.005 13.700 4.235 ;
        RECT  10.430 3.010 10.470 4.235 ;
        RECT  10.420 2.710 10.430 4.235 ;
        RECT  10.345 2.660 10.420 4.235 ;
        RECT  10.240 2.405 10.345 4.235 ;
        RECT  10.115 2.405 10.240 3.240 ;
        RECT  10.090 2.630 10.115 3.240 ;
        RECT  9.510 3.010 10.090 3.240 ;
        RECT  9.280 3.010 9.510 4.405 ;
        RECT  6.820 4.175 9.280 4.405 ;
        RECT  6.590 3.445 6.820 4.405 ;
        RECT  5.895 3.445 6.590 3.675 ;
        RECT  5.665 3.445 5.895 4.410 ;
        RECT  3.990 4.180 5.665 4.410 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.575 2.250 13.315 2.690 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.600 1.845 15.625 2.075 ;
        RECT  15.370 1.330 15.600 3.610 ;
        RECT  14.560 1.330 15.370 1.560 ;
        RECT  15.005 3.380 15.370 3.610 ;
        RECT  14.665 3.380 15.005 3.720 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.850 2.060 1.400 2.765 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 3.810 0.625 4.150 ;
        RECT  0.150 3.810 0.620 4.390 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.450 -0.400 15.840 0.400 ;
        RECT  13.110 -0.400 13.450 1.555 ;
        RECT  9.790 -0.400 13.110 0.400 ;
        RECT  9.450 -0.400 9.790 0.575 ;
        RECT  7.110 -0.400 9.450 0.400 ;
        RECT  6.770 -0.400 7.110 1.075 ;
        RECT  3.665 -0.400 6.770 0.400 ;
        RECT  3.325 -0.400 3.665 0.900 ;
        RECT  1.205 -0.400 3.325 0.400 ;
        RECT  0.865 -0.400 1.205 0.575 ;
        RECT  0.000 -0.400 0.865 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.660 4.640 15.840 5.440 ;
        RECT  15.320 4.465 15.660 5.440 ;
        RECT  13.655 4.640 15.320 5.440 ;
        RECT  13.315 4.465 13.655 5.440 ;
        RECT  12.345 4.640 13.315 5.440 ;
        RECT  12.005 4.465 12.345 5.440 ;
        RECT  10.010 4.640 12.005 5.440 ;
        RECT  9.780 3.640 10.010 5.440 ;
        RECT  6.355 4.640 9.780 5.440 ;
        RECT  6.125 3.915 6.355 5.440 ;
        RECT  3.660 4.640 6.125 5.440 ;
        RECT  3.320 4.465 3.660 5.440 ;
        RECT  1.195 4.640 3.320 5.440 ;
        RECT  0.855 4.465 1.195 5.440 ;
        RECT  0.000 4.640 0.855 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.510 0.870 15.660 1.100 ;
        RECT  15.280 0.795 15.510 1.100 ;
        RECT  14.205 0.795 15.280 1.025 ;
        RECT  14.980 1.940 15.090 2.280 ;
        RECT  14.750 1.790 14.980 2.280 ;
        RECT  12.690 1.790 14.750 2.020 ;
        RECT  14.170 0.795 14.205 1.500 ;
        RECT  13.975 0.795 14.170 1.555 ;
        RECT  13.830 1.215 13.975 1.555 ;
        RECT  13.210 2.975 13.320 3.205 ;
        RECT  12.980 2.975 13.210 3.775 ;
        RECT  12.345 2.975 12.980 3.205 ;
        RECT  11.885 3.545 12.980 3.775 ;
        RECT  12.350 1.420 12.690 2.020 ;
        RECT  12.345 1.790 12.350 2.020 ;
        RECT  12.115 1.790 12.345 3.205 ;
        RECT  12.000 0.720 12.190 1.060 ;
        RECT  11.850 0.720 12.000 1.505 ;
        RECT  11.655 2.480 11.885 3.775 ;
        RECT  11.770 0.775 11.850 1.505 ;
        RECT  10.250 1.275 11.770 1.505 ;
        RECT  11.335 1.740 11.390 1.970 ;
        RECT  10.930 1.735 11.335 1.980 ;
        RECT  11.005 0.660 11.060 1.000 ;
        RECT  10.720 0.660 11.005 1.035 ;
        RECT  10.700 1.735 10.930 3.580 ;
        RECT  9.910 0.805 10.720 1.035 ;
        RECT  9.530 1.750 10.700 2.015 ;
        RECT  9.680 0.805 9.910 1.270 ;
        RECT  9.045 1.040 9.680 1.270 ;
        RECT  9.295 1.750 9.530 2.120 ;
        RECT  8.815 1.040 9.045 3.225 ;
        RECT  8.645 3.605 8.985 3.945 ;
        RECT  8.290 1.040 8.815 1.270 ;
        RECT  8.220 2.995 8.815 3.225 ;
        RECT  7.280 3.715 8.645 3.945 ;
        RECT  8.350 1.500 8.580 2.710 ;
        RECT  7.870 1.500 8.350 1.730 ;
        RECT  7.740 2.480 8.350 2.710 ;
        RECT  7.280 1.960 8.110 2.190 ;
        RECT  7.640 1.070 7.870 1.730 ;
        RECT  7.510 2.480 7.740 3.480 ;
        RECT  7.530 1.070 7.640 1.410 ;
        RECT  7.050 1.310 7.280 3.945 ;
        RECT  6.310 1.310 7.050 1.540 ;
        RECT  6.050 2.975 7.050 3.205 ;
        RECT  6.465 2.255 6.780 2.485 ;
        RECT  6.235 1.775 6.465 2.485 ;
        RECT  6.150 1.200 6.310 1.540 ;
        RECT  5.005 1.775 6.235 2.005 ;
        RECT  5.970 0.630 6.150 1.540 ;
        RECT  5.920 0.630 5.970 1.485 ;
        RECT  5.615 2.240 5.955 2.580 ;
        RECT  5.810 0.630 5.920 0.970 ;
        RECT  5.430 2.350 5.615 2.580 ;
        RECT  5.200 2.350 5.430 3.845 ;
        RECT  2.840 3.615 5.200 3.845 ;
        RECT  4.970 1.300 5.005 2.005 ;
        RECT  4.740 1.300 4.970 3.270 ;
        RECT  4.665 1.300 4.740 1.640 ;
        RECT  4.320 3.040 4.740 3.270 ;
        RECT  4.280 2.005 4.510 2.380 ;
        RECT  3.980 3.040 4.320 3.380 ;
        RECT  2.625 2.005 4.280 2.235 ;
        RECT  3.400 3.040 3.980 3.270 ;
        RECT  3.390 2.525 3.400 3.270 ;
        RECT  3.170 2.470 3.390 3.270 ;
        RECT  3.050 2.470 3.170 2.810 ;
        RECT  2.610 3.615 2.840 4.345 ;
        RECT  2.395 1.195 2.625 2.735 ;
        RECT  1.885 4.115 2.610 4.345 ;
        RECT  2.100 1.195 2.395 1.425 ;
        RECT  2.345 2.505 2.395 2.735 ;
        RECT  2.115 2.505 2.345 3.825 ;
        RECT  1.885 1.770 2.150 2.110 ;
        RECT  1.810 1.770 1.885 4.345 ;
        RECT  1.655 1.825 1.810 4.345 ;
        RECT  0.520 3.220 1.655 3.450 ;
        RECT  0.465 1.210 0.520 1.550 ;
        RECT  0.465 3.165 0.520 3.505 ;
        RECT  0.235 1.210 0.465 3.505 ;
        RECT  0.180 1.210 0.235 1.550 ;
        RECT  0.180 3.165 0.235 3.505 ;
    END
END DFFSRHQX1

MACRO DFFSRXL
    CLASS CORE ;
    FOREIGN DFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.360 4.035 11.730 4.365 ;
        RECT  8.795 4.135 11.360 4.365 ;
        RECT  8.490 4.125 8.795 4.365 ;
        RECT  6.155 4.125 8.490 4.355 ;
        RECT  6.095 4.085 6.155 4.355 ;
        RECT  5.865 4.005 6.095 4.355 ;
        RECT  5.040 4.005 5.865 4.235 ;
        RECT  4.810 4.005 5.040 4.365 ;
        RECT  4.540 4.135 4.810 4.365 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.625 1.790 6.680 2.130 ;
        RECT  6.155 1.785 6.625 2.175 ;
        RECT  6.075 1.785 6.155 2.155 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.120 1.095 15.360 1.435 ;
        RECT  14.890 1.095 15.120 3.455 ;
        RECT  14.715 2.965 14.890 3.455 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.555 1.095 16.685 1.435 ;
        RECT  16.345 1.095 16.555 3.230 ;
        RECT  16.330 1.205 16.345 3.230 ;
        RECT  16.325 1.205 16.330 3.580 ;
        RECT  15.990 2.965 16.325 3.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.215 2.155 0.875 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  8.010 2.250 8.575 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.125 -0.400 17.160 0.400 ;
        RECT  15.785 -0.400 16.125 0.575 ;
        RECT  14.650 -0.400 15.785 0.400 ;
        RECT  14.310 -0.400 14.650 0.575 ;
        RECT  11.455 -0.400 14.310 0.400 ;
        RECT  11.115 -0.400 11.455 0.575 ;
        RECT  8.890 -0.400 11.115 0.400 ;
        RECT  8.550 -0.400 8.890 1.485 ;
        RECT  7.115 -0.400 8.550 0.400 ;
        RECT  6.885 -0.400 7.115 0.900 ;
        RECT  4.195 -0.400 6.885 0.400 ;
        RECT  3.855 -0.400 4.195 0.900 ;
        RECT  1.330 -0.400 3.855 0.400 ;
        RECT  0.990 -0.400 1.330 0.575 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.095 4.640 17.160 5.440 ;
        RECT  15.720 4.465 16.095 5.440 ;
        RECT  13.570 4.640 15.720 5.440 ;
        RECT  13.230 3.395 13.570 5.440 ;
        RECT  12.405 4.640 13.230 5.440 ;
        RECT  12.175 3.395 12.405 5.440 ;
        RECT  11.490 3.395 12.175 3.625 ;
        RECT  5.635 4.640 12.175 5.440 ;
        RECT  11.130 3.310 11.490 3.625 ;
        RECT  10.905 3.395 11.130 3.625 ;
        RECT  10.675 3.395 10.905 3.845 ;
        RECT  8.795 3.615 10.675 3.845 ;
        RECT  8.510 3.460 8.795 3.845 ;
        RECT  8.455 3.460 8.510 3.800 ;
        RECT  5.295 4.465 5.635 5.440 ;
        RECT  4.310 4.640 5.295 5.440 ;
        RECT  3.970 4.465 4.310 5.440 ;
        RECT  1.340 4.640 3.970 5.440 ;
        RECT  0.945 4.465 1.340 5.440 ;
        RECT  0.000 4.640 0.945 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.600 2.220 15.920 2.560 ;
        RECT  15.580 2.220 15.600 3.915 ;
        RECT  15.370 2.275 15.580 3.915 ;
        RECT  14.475 3.685 15.370 3.915 ;
        RECT  14.415 1.170 14.660 1.510 ;
        RECT  14.415 3.505 14.475 3.915 ;
        RECT  14.320 1.170 14.415 3.915 ;
        RECT  14.245 1.225 14.320 3.915 ;
        RECT  14.185 1.225 14.245 3.735 ;
        RECT  13.950 3.395 14.185 3.735 ;
        RECT  13.725 1.825 13.955 3.165 ;
        RECT  13.605 0.980 13.855 1.320 ;
        RECT  13.145 1.825 13.725 2.055 ;
        RECT  12.010 2.935 13.725 3.165 ;
        RECT  13.515 0.630 13.605 1.320 ;
        RECT  13.375 0.630 13.515 1.265 ;
        RECT  12.275 0.630 13.375 0.860 ;
        RECT  12.915 1.090 13.145 2.055 ;
        RECT  12.715 1.090 12.915 1.320 ;
        RECT  12.135 1.890 12.475 2.230 ;
        RECT  12.255 0.630 12.275 1.235 ;
        RECT  12.045 0.630 12.255 1.290 ;
        RECT  11.065 1.890 12.135 2.120 ;
        RECT  11.915 0.950 12.045 1.290 ;
        RECT  11.780 2.615 12.010 3.165 ;
        RECT  11.295 2.615 11.780 2.845 ;
        RECT  10.955 2.560 11.295 2.900 ;
        RECT  10.835 1.250 11.065 2.120 ;
        RECT  10.415 1.250 10.835 1.480 ;
        RECT  9.545 0.720 10.705 0.950 ;
        RECT  10.185 1.250 10.415 3.360 ;
        RECT  10.115 1.250 10.185 1.535 ;
        RECT  9.775 3.130 10.185 3.360 ;
        RECT  9.885 1.195 10.115 1.535 ;
        RECT  9.545 2.430 9.870 2.770 ;
        RECT  9.315 0.720 9.545 3.125 ;
        RECT  8.035 1.745 9.315 1.975 ;
        RECT  8.075 2.895 9.315 3.125 ;
        RECT  8.020 2.895 8.075 3.800 ;
        RECT  7.805 1.370 8.035 1.975 ;
        RECT  7.845 2.895 8.020 3.835 ;
        RECT  7.575 0.740 7.935 0.970 ;
        RECT  7.735 3.460 7.845 3.835 ;
        RECT  6.555 3.605 7.735 3.835 ;
        RECT  7.345 0.740 7.575 1.365 ;
        RECT  5.670 1.135 7.345 1.365 ;
        RECT  7.260 1.635 7.300 2.795 ;
        RECT  7.245 1.635 7.260 2.800 ;
        RECT  7.070 1.635 7.245 3.375 ;
        RECT  6.920 2.460 7.070 3.375 ;
        RECT  6.870 2.565 6.920 3.375 ;
        RECT  6.785 2.905 6.870 3.375 ;
        RECT  6.100 2.905 6.785 3.135 ;
        RECT  6.325 3.545 6.555 3.835 ;
        RECT  3.720 3.545 6.325 3.775 ;
        RECT  5.870 2.540 6.100 3.135 ;
        RECT  5.640 1.120 5.670 1.460 ;
        RECT  5.410 1.120 5.640 3.135 ;
        RECT  5.330 1.120 5.410 1.460 ;
        RECT  5.090 2.905 5.410 3.135 ;
        RECT  4.935 1.840 5.165 2.205 ;
        RECT  4.045 2.905 5.090 3.260 ;
        RECT  3.585 1.975 4.935 2.205 ;
        RECT  3.815 2.510 4.045 3.260 ;
        RECT  3.490 3.545 3.720 4.365 ;
        RECT  3.355 0.955 3.585 2.965 ;
        RECT  3.140 4.135 3.490 4.365 ;
        RECT  3.030 0.955 3.355 1.240 ;
        RECT  3.055 2.735 3.355 2.965 ;
        RECT  2.895 1.770 3.125 2.225 ;
        RECT  3.055 3.480 3.110 3.820 ;
        RECT  2.825 2.735 3.055 3.820 ;
        RECT  2.690 0.900 3.030 1.240 ;
        RECT  2.430 1.995 2.895 2.225 ;
        RECT  2.770 3.480 2.825 3.820 ;
        RECT  2.430 3.045 2.505 3.405 ;
        RECT  2.230 1.490 2.430 3.405 ;
        RECT  2.275 3.980 2.330 4.320 ;
        RECT  1.990 3.810 2.275 4.320 ;
        RECT  2.215 1.435 2.230 3.405 ;
        RECT  1.845 0.745 2.225 1.050 ;
        RECT  2.200 1.435 2.215 3.300 ;
        RECT  1.890 1.435 2.200 1.775 ;
        RECT  1.555 2.960 2.200 3.300 ;
        RECT  0.520 3.810 1.990 4.040 ;
        RECT  0.465 0.815 1.845 1.045 ;
        RECT  0.465 1.430 0.520 1.770 ;
        RECT  0.290 3.000 0.520 4.040 ;
        RECT  0.235 0.815 0.465 1.770 ;
        RECT  0.180 3.000 0.290 3.340 ;
        RECT  0.180 1.430 0.235 1.770 ;
    END
END DFFSRXL

MACRO DFFSRX4
    CLASS CORE ;
    FOREIGN DFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRXL ;
    SIZE 23.760 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.180 3.995 14.520 4.335 ;
        RECT  9.025 4.000 14.180 4.230 ;
        RECT  8.700 4.000 9.025 4.335 ;
        RECT  4.860 4.105 8.700 4.335 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.795 2.295 7.265 2.790 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.565 1.820 21.640 3.220 ;
        RECT  21.335 1.475 21.565 3.220 ;
        RECT  21.260 1.420 21.335 3.220 ;
        RECT  21.255 1.420 21.260 3.195 ;
        RECT  20.860 1.420 21.255 1.820 ;
        RECT  20.900 2.855 21.255 3.195 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.885 1.820 22.960 3.220 ;
        RECT  22.655 1.475 22.885 3.220 ;
        RECT  22.580 1.420 22.655 3.220 ;
        RECT  22.240 1.420 22.580 1.860 ;
        RECT  22.265 2.855 22.580 3.195 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 2.445 0.930 2.785 ;
        RECT  0.140 2.405 0.730 2.785 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.510 2.385 1.620 2.725 ;
        RECT  1.280 1.870 1.510 2.725 ;
        RECT  1.105 1.870 1.280 2.100 ;
        RECT  0.875 1.845 1.105 2.100 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.260 -0.400 23.760 0.400 ;
        RECT  22.920 -0.400 23.260 0.575 ;
        RECT  21.880 -0.400 22.920 0.400 ;
        RECT  21.540 -0.400 21.880 0.575 ;
        RECT  20.520 -0.400 21.540 0.400 ;
        RECT  20.180 -0.400 20.520 0.575 ;
        RECT  15.350 -0.400 20.180 0.400 ;
        RECT  15.010 -0.400 15.350 1.050 ;
        RECT  12.465 -0.400 15.010 0.400 ;
        RECT  12.125 -0.400 12.465 1.145 ;
        RECT  9.865 -0.400 12.125 0.400 ;
        RECT  9.525 -0.400 9.865 1.320 ;
        RECT  7.260 -0.400 9.525 0.400 ;
        RECT  6.920 -0.400 7.260 0.860 ;
        RECT  4.540 -0.400 6.920 0.400 ;
        RECT  4.200 -0.400 4.540 0.845 ;
        RECT  1.295 -0.400 4.200 0.400 ;
        RECT  0.955 -0.400 1.295 0.575 ;
        RECT  0.000 -0.400 0.955 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.285 4.640 23.760 5.440 ;
        RECT  22.945 4.465 23.285 5.440 ;
        RECT  21.920 4.640 22.945 5.440 ;
        RECT  21.580 4.465 21.920 5.440 ;
        RECT  20.560 4.640 21.580 5.440 ;
        RECT  20.220 4.465 20.560 5.440 ;
        RECT  17.810 4.640 20.220 5.440 ;
        RECT  17.470 3.640 17.810 5.440 ;
        RECT  15.805 4.640 17.470 5.440 ;
        RECT  15.465 2.920 15.805 5.440 ;
        RECT  13.545 4.640 15.465 5.440 ;
        RECT  13.205 4.465 13.545 5.440 ;
        RECT  12.390 4.640 13.205 5.440 ;
        RECT  12.050 4.465 12.390 5.440 ;
        RECT  9.725 4.640 12.050 5.440 ;
        RECT  9.385 4.465 9.725 5.440 ;
        RECT  4.610 4.640 9.385 5.440 ;
        RECT  4.270 4.465 4.610 5.440 ;
        RECT  1.095 4.640 4.270 5.440 ;
        RECT  0.755 4.465 1.095 5.440 ;
        RECT  0.000 4.640 0.755 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  23.195 2.210 23.425 3.740 ;
        RECT  20.495 3.510 23.195 3.740 ;
        RECT  20.265 1.670 20.495 3.740 ;
        RECT  19.700 1.670 20.265 1.900 ;
        RECT  19.800 3.400 20.265 3.740 ;
        RECT  19.240 2.160 19.950 2.500 ;
        RECT  19.460 3.260 19.800 4.070 ;
        RECT  19.470 0.920 19.700 1.900 ;
        RECT  19.100 1.375 19.240 3.015 ;
        RECT  19.010 1.375 19.100 3.845 ;
        RECT  18.250 1.375 19.010 1.605 ;
        RECT  18.870 2.785 19.010 3.845 ;
        RECT  18.685 0.675 18.915 1.030 ;
        RECT  18.760 3.035 18.870 3.845 ;
        RECT  18.720 1.920 18.775 2.260 ;
        RECT  16.530 3.085 18.760 3.315 ;
        RECT  18.435 1.860 18.720 2.260 ;
        RECT  17.530 0.675 18.685 0.905 ;
        RECT  16.310 1.860 18.435 2.090 ;
        RECT  17.880 1.205 18.250 1.605 ;
        RECT  16.905 1.375 17.880 1.605 ;
        RECT  17.190 0.675 17.530 1.050 ;
        RECT  16.075 0.675 17.190 0.905 ;
        RECT  16.675 1.140 16.905 1.605 ;
        RECT  16.465 1.140 16.675 1.370 ;
        RECT  16.420 3.025 16.530 3.835 ;
        RECT  16.190 2.455 16.420 3.835 ;
        RECT  16.025 1.860 16.310 2.155 ;
        RECT  15.085 2.455 16.190 2.685 ;
        RECT  15.965 0.675 16.075 1.290 ;
        RECT  13.880 1.925 16.025 2.155 ;
        RECT  15.845 0.675 15.965 1.605 ;
        RECT  15.735 0.950 15.845 1.605 ;
        RECT  14.630 1.375 15.735 1.605 ;
        RECT  15.130 4.070 15.235 4.410 ;
        RECT  14.900 3.535 15.130 4.410 ;
        RECT  15.030 2.455 15.085 3.150 ;
        RECT  14.855 2.455 15.030 3.305 ;
        RECT  8.395 3.535 14.900 3.765 ;
        RECT  14.895 4.070 14.900 4.410 ;
        RECT  14.745 2.810 14.855 3.305 ;
        RECT  12.955 3.075 14.745 3.305 ;
        RECT  14.400 0.970 14.630 1.605 ;
        RECT  14.290 0.970 14.400 1.310 ;
        RECT  13.650 0.880 13.880 2.155 ;
        RECT  13.485 0.880 13.650 1.110 ;
        RECT  13.490 1.925 13.650 2.155 ;
        RECT  13.260 1.925 13.490 2.845 ;
        RECT  13.080 1.355 13.420 1.695 ;
        RECT  11.255 1.925 13.260 2.155 ;
        RECT  11.720 1.410 13.080 1.640 ;
        RECT  12.725 2.385 12.955 3.305 ;
        RECT  12.520 2.385 12.725 2.615 ;
        RECT  11.490 0.675 11.720 1.640 ;
        RECT  10.455 0.675 11.490 0.905 ;
        RECT  11.145 1.755 11.255 3.135 ;
        RECT  11.055 1.220 11.145 3.135 ;
        RECT  11.025 1.220 11.055 3.190 ;
        RECT  10.915 1.220 11.025 1.985 ;
        RECT  10.715 2.850 11.025 3.190 ;
        RECT  10.805 1.220 10.915 1.560 ;
        RECT  10.455 2.245 10.790 2.585 ;
        RECT  10.450 0.675 10.455 2.585 ;
        RECT  10.225 0.675 10.450 2.530 ;
        RECT  8.895 2.045 10.225 2.275 ;
        RECT  8.765 1.400 9.105 1.740 ;
        RECT  8.860 2.910 9.105 3.250 ;
        RECT  7.765 0.745 8.915 0.975 ;
        RECT  8.765 2.565 8.860 3.250 ;
        RECT  8.600 1.455 8.765 1.740 ;
        RECT  8.630 2.565 8.765 3.195 ;
        RECT  8.600 2.565 8.630 2.795 ;
        RECT  8.370 1.455 8.600 2.795 ;
        RECT  8.165 3.085 8.395 3.765 ;
        RECT  8.145 2.220 8.370 2.450 ;
        RECT  7.805 3.085 8.165 3.315 ;
        RECT  7.805 1.625 7.955 1.855 ;
        RECT  7.880 3.605 7.935 3.835 ;
        RECT  7.650 3.605 7.880 3.840 ;
        RECT  7.575 1.625 7.805 3.315 ;
        RECT  7.535 0.745 7.765 1.345 ;
        RECT  3.885 3.610 7.650 3.840 ;
        RECT  6.370 3.085 7.575 3.315 ;
        RECT  5.900 1.115 7.535 1.345 ;
        RECT  6.140 2.280 6.370 3.315 ;
        RECT  5.670 1.115 5.900 3.375 ;
        RECT  5.600 1.115 5.670 1.435 ;
        RECT  4.265 3.145 5.670 3.375 ;
        RECT  5.205 1.775 5.435 2.240 ;
        RECT  3.425 1.775 5.205 2.005 ;
        RECT  4.265 2.330 4.320 2.670 ;
        RECT  4.035 2.330 4.265 3.375 ;
        RECT  3.980 2.330 4.035 2.670 ;
        RECT  3.655 3.610 3.885 4.410 ;
        RECT  2.790 4.180 3.655 4.410 ;
        RECT  3.355 0.665 3.425 2.005 ;
        RECT  3.250 0.665 3.355 2.415 ;
        RECT  3.125 0.665 3.250 3.805 ;
        RECT  3.040 0.665 3.125 0.895 ;
        RECT  3.020 2.185 3.125 3.805 ;
        RECT  2.175 1.520 2.810 1.860 ;
        RECT  2.560 3.130 2.790 4.410 ;
        RECT  2.275 0.630 2.655 1.045 ;
        RECT  2.175 3.130 2.560 3.360 ;
        RECT  2.030 3.740 2.330 4.100 ;
        RECT  0.735 0.815 2.275 1.045 ;
        RECT  1.945 1.445 2.175 3.360 ;
        RECT  0.520 3.815 2.030 4.045 ;
        RECT  1.765 1.445 1.945 1.675 ;
        RECT  1.505 3.020 1.945 3.360 ;
        RECT  0.505 0.815 0.735 1.555 ;
        RECT  0.290 3.215 0.520 4.045 ;
        RECT  0.395 1.325 0.505 1.555 ;
        RECT  0.180 3.215 0.290 3.555 ;
    END
END DFFSRX4

MACRO DFFSRX2
    CLASS CORE ;
    FOREIGN DFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.170 4.035 11.665 4.365 ;
        RECT  11.005 4.085 11.170 4.365 ;
        RECT  8.525 4.135 11.005 4.365 ;
        RECT  8.295 4.125 8.525 4.365 ;
        RECT  5.900 4.125 8.295 4.355 ;
        RECT  5.670 4.005 5.900 4.355 ;
        RECT  4.845 4.005 5.670 4.235 ;
        RECT  4.615 4.005 4.845 4.365 ;
        RECT  4.345 4.135 4.615 4.365 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.085 1.770 6.625 2.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.140 1.190 15.295 1.530 ;
        RECT  14.965 1.190 15.140 3.205 ;
        RECT  14.910 1.190 14.965 3.335 ;
        RECT  14.680 2.965 14.910 3.335 ;
        RECT  14.625 3.105 14.680 3.335 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.840 2.955 16.945 3.195 ;
        RECT  16.820 1.105 16.840 3.195 ;
        RECT  16.815 1.105 16.820 4.140 ;
        RECT  16.610 1.050 16.815 4.140 ;
        RECT  16.475 1.050 16.610 1.390 ;
        RECT  16.560 2.965 16.610 4.140 ;
        RECT  16.355 3.200 16.560 4.140 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.565 2.115 1.180 2.730 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  7.815 2.250 8.605 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.055 -0.400 17.160 0.400 ;
        RECT  15.715 -0.400 16.055 1.690 ;
        RECT  14.320 -0.400 15.715 0.400 ;
        RECT  13.980 -0.400 14.320 0.575 ;
        RECT  11.280 -0.400 13.980 0.400 ;
        RECT  10.940 -0.400 11.280 0.575 ;
        RECT  8.695 -0.400 10.940 0.400 ;
        RECT  8.355 -0.400 8.695 1.400 ;
        RECT  6.960 -0.400 8.355 0.400 ;
        RECT  6.730 -0.400 6.960 0.900 ;
        RECT  4.000 -0.400 6.730 0.400 ;
        RECT  3.660 -0.400 4.000 0.900 ;
        RECT  1.335 -0.400 3.660 0.400 ;
        RECT  0.995 -0.400 1.335 0.575 ;
        RECT  0.000 -0.400 0.995 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.875 4.640 17.160 5.440 ;
        RECT  15.535 4.090 15.875 5.440 ;
        RECT  13.295 4.640 15.535 5.440 ;
        RECT  12.955 3.560 13.295 5.440 ;
        RECT  12.210 4.640 12.955 5.440 ;
        RECT  11.980 3.485 12.210 5.440 ;
        RECT  10.710 3.485 11.980 3.715 ;
        RECT  5.440 4.640 11.980 5.440 ;
        RECT  10.480 3.485 10.710 3.845 ;
        RECT  8.640 3.615 10.480 3.845 ;
        RECT  8.300 3.505 8.640 3.845 ;
        RECT  5.100 4.465 5.440 5.440 ;
        RECT  4.115 4.640 5.100 5.440 ;
        RECT  3.775 4.465 4.115 5.440 ;
        RECT  1.280 4.640 3.775 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.750 2.145 16.255 2.375 ;
        RECT  15.520 2.145 15.750 3.830 ;
        RECT  14.380 3.600 15.520 3.830 ;
        RECT  14.340 1.225 14.380 3.950 ;
        RECT  14.150 1.170 14.340 3.950 ;
        RECT  14.000 1.170 14.150 1.510 ;
        RECT  14.020 3.665 14.150 3.950 ;
        RECT  13.680 3.665 14.020 4.005 ;
        RECT  13.610 1.825 13.840 3.165 ;
        RECT  12.825 1.825 13.610 2.055 ;
        RECT  12.015 2.935 13.610 3.165 ;
        RECT  13.465 0.780 13.520 1.120 ;
        RECT  13.180 0.745 13.465 1.120 ;
        RECT  12.080 0.745 13.180 0.975 ;
        RECT  12.595 1.275 12.825 2.055 ;
        RECT  12.460 1.275 12.595 1.505 ;
        RECT  11.995 1.855 12.225 2.230 ;
        RECT  11.795 0.745 12.080 1.120 ;
        RECT  11.675 2.880 12.015 3.220 ;
        RECT  10.870 1.855 11.995 2.085 ;
        RECT  11.740 0.780 11.795 1.120 ;
        RECT  11.620 2.880 11.675 3.110 ;
        RECT  11.390 2.615 11.620 3.110 ;
        RECT  10.535 2.615 11.390 2.845 ;
        RECT  10.640 1.335 10.870 2.085 ;
        RECT  10.220 1.335 10.640 1.565 ;
        RECT  9.345 0.735 10.510 0.965 ;
        RECT  9.990 1.335 10.220 3.270 ;
        RECT  9.975 1.335 9.990 1.620 ;
        RECT  9.920 3.040 9.990 3.270 ;
        RECT  9.635 1.280 9.975 1.620 ;
        RECT  9.580 3.040 9.920 3.380 ;
        RECT  9.365 2.525 9.675 2.755 ;
        RECT  9.345 1.745 9.365 2.755 ;
        RECT  9.115 0.735 9.345 3.225 ;
        RECT  7.880 1.745 9.115 1.975 ;
        RECT  7.920 2.995 9.115 3.225 ;
        RECT  7.690 2.995 7.920 3.835 ;
        RECT  7.650 1.370 7.880 1.975 ;
        RECT  7.420 0.745 7.740 0.975 ;
        RECT  7.580 3.460 7.690 3.835 ;
        RECT  6.360 3.605 7.580 3.835 ;
        RECT  7.190 0.745 7.420 1.365 ;
        RECT  7.110 2.460 7.200 2.800 ;
        RECT  5.475 1.135 7.190 1.365 ;
        RECT  6.880 1.600 7.110 3.375 ;
        RECT  6.860 2.460 6.880 3.375 ;
        RECT  6.820 2.515 6.860 3.375 ;
        RECT  6.590 2.905 6.820 3.375 ;
        RECT  5.905 2.905 6.590 3.135 ;
        RECT  6.130 3.545 6.360 3.835 ;
        RECT  3.525 3.545 6.130 3.775 ;
        RECT  5.675 2.540 5.905 3.135 ;
        RECT  5.445 1.120 5.475 1.460 ;
        RECT  5.215 1.120 5.445 3.135 ;
        RECT  5.135 1.120 5.215 1.460 ;
        RECT  4.895 2.905 5.215 3.135 ;
        RECT  4.740 1.840 4.970 2.205 ;
        RECT  3.850 2.905 4.895 3.260 ;
        RECT  3.390 1.975 4.740 2.205 ;
        RECT  3.620 2.510 3.850 3.260 ;
        RECT  3.295 3.545 3.525 4.365 ;
        RECT  3.160 0.955 3.390 2.965 ;
        RECT  2.945 4.135 3.295 4.365 ;
        RECT  2.835 0.955 3.160 1.240 ;
        RECT  2.860 2.735 3.160 2.965 ;
        RECT  2.700 1.770 2.930 2.225 ;
        RECT  2.630 2.735 2.860 3.820 ;
        RECT  2.495 0.900 2.835 1.240 ;
        RECT  2.235 1.995 2.700 2.225 ;
        RECT  2.235 3.180 2.330 3.655 ;
        RECT  2.035 1.455 2.235 3.655 ;
        RECT  1.810 3.980 2.150 4.320 ;
        RECT  1.660 0.695 2.070 1.060 ;
        RECT  2.005 1.400 2.035 3.655 ;
        RECT  1.695 1.400 2.005 1.740 ;
        RECT  1.500 3.180 2.005 3.465 ;
        RECT  0.520 3.980 1.810 4.210 ;
        RECT  0.640 0.830 1.660 1.060 ;
        RECT  0.635 0.830 0.640 1.625 ;
        RECT  0.410 0.830 0.635 1.680 ;
        RECT  0.290 3.150 0.520 4.210 ;
        RECT  0.295 1.340 0.410 1.680 ;
        RECT  0.180 3.150 0.290 3.490 ;
    END
END DFFSRX2

MACRO DFFSRX1
    CLASS CORE ;
    FOREIGN DFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 4.035 11.725 4.265 ;
        RECT  11.360 4.035 11.665 4.365 ;
        RECT  8.795 4.135 11.360 4.365 ;
        RECT  8.485 4.125 8.795 4.365 ;
        RECT  6.155 4.125 8.485 4.355 ;
        RECT  6.090 4.085 6.155 4.355 ;
        RECT  5.860 4.005 6.090 4.355 ;
        RECT  5.035 4.005 5.860 4.235 ;
        RECT  4.805 4.005 5.035 4.365 ;
        RECT  4.535 4.135 4.805 4.365 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.080 1.765 6.620 2.230 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.115 1.155 15.230 1.495 ;
        RECT  15.115 3.115 15.155 3.455 ;
        RECT  14.890 1.155 15.115 3.455 ;
        RECT  14.885 1.165 14.890 3.455 ;
        RECT  14.815 2.965 14.885 3.455 ;
        RECT  14.735 2.965 14.815 3.400 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.550 1.245 16.650 3.185 ;
        RECT  16.475 1.190 16.550 3.185 ;
        RECT  16.420 1.190 16.475 3.730 ;
        RECT  16.285 1.190 16.420 1.540 ;
        RECT  16.360 2.940 16.420 3.730 ;
        RECT  16.135 2.955 16.360 3.730 ;
        RECT  16.210 1.190 16.285 1.530 ;
        RECT  16.130 2.955 16.135 3.725 ;
        RECT  16.055 2.955 16.130 3.195 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.280 1.400 2.660 ;
        RECT  0.635 2.280 0.800 2.620 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  8.005 2.250 8.580 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.865 -0.400 17.160 0.400 ;
        RECT  15.525 -0.400 15.865 0.575 ;
        RECT  14.510 -0.400 15.525 0.400 ;
        RECT  14.170 -0.400 14.510 0.575 ;
        RECT  11.470 -0.400 14.170 0.400 ;
        RECT  11.130 -0.400 11.470 0.575 ;
        RECT  8.885 -0.400 11.130 0.400 ;
        RECT  8.545 -0.400 8.885 1.485 ;
        RECT  7.110 -0.400 8.545 0.400 ;
        RECT  6.880 -0.400 7.110 0.900 ;
        RECT  4.190 -0.400 6.880 0.400 ;
        RECT  3.850 -0.400 4.190 0.900 ;
        RECT  1.425 -0.400 3.850 0.400 ;
        RECT  1.085 -0.400 1.425 0.575 ;
        RECT  0.000 -0.400 1.085 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.760 4.640 17.160 5.440 ;
        RECT  15.420 4.465 15.760 5.440 ;
        RECT  13.565 4.640 15.420 5.440 ;
        RECT  13.225 3.395 13.565 5.440 ;
        RECT  12.400 4.640 13.225 5.440 ;
        RECT  12.170 3.430 12.400 5.440 ;
        RECT  10.900 3.430 12.170 3.660 ;
        RECT  5.630 4.640 12.170 5.440 ;
        RECT  10.670 3.430 10.900 3.845 ;
        RECT  8.960 3.615 10.670 3.845 ;
        RECT  8.790 3.455 8.960 3.845 ;
        RECT  8.730 3.400 8.790 3.845 ;
        RECT  8.450 3.400 8.730 3.740 ;
        RECT  5.290 4.465 5.630 5.440 ;
        RECT  4.305 4.640 5.290 5.440 ;
        RECT  3.965 4.465 4.305 5.440 ;
        RECT  1.130 4.640 3.965 5.440 ;
        RECT  0.790 4.465 1.130 5.440 ;
        RECT  0.000 4.640 0.790 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.740 2.210 16.080 2.550 ;
        RECT  15.620 2.320 15.740 2.550 ;
        RECT  15.390 2.320 15.620 4.040 ;
        RECT  14.310 3.810 15.390 4.040 ;
        RECT  14.310 1.170 14.530 1.510 ;
        RECT  14.190 1.170 14.310 4.040 ;
        RECT  14.080 1.225 14.190 4.040 ;
        RECT  13.945 3.395 14.080 3.735 ;
        RECT  13.605 2.110 13.715 2.450 ;
        RECT  13.600 0.980 13.710 1.320 ;
        RECT  13.375 1.825 13.605 3.165 ;
        RECT  13.370 0.630 13.600 1.320 ;
        RECT  13.015 1.825 13.375 2.055 ;
        RECT  11.810 2.935 13.375 3.165 ;
        RECT  12.270 0.630 13.370 0.860 ;
        RECT  12.785 1.090 13.015 2.055 ;
        RECT  12.650 1.090 12.785 1.320 ;
        RECT  12.185 1.855 12.415 2.230 ;
        RECT  12.040 0.630 12.270 1.290 ;
        RECT  11.060 1.855 12.185 2.085 ;
        RECT  11.930 0.950 12.040 1.290 ;
        RECT  11.580 2.615 11.810 3.165 ;
        RECT  10.725 2.615 11.580 2.845 ;
        RECT  10.830 1.250 11.060 2.085 ;
        RECT  10.410 1.250 10.830 1.480 ;
        RECT  9.535 0.735 10.700 0.965 ;
        RECT  10.180 1.250 10.410 3.330 ;
        RECT  10.165 1.250 10.180 1.535 ;
        RECT  9.770 3.100 10.180 3.330 ;
        RECT  9.825 1.195 10.165 1.535 ;
        RECT  9.555 2.525 9.865 2.755 ;
        RECT  9.535 1.745 9.555 2.755 ;
        RECT  9.305 0.735 9.535 3.125 ;
        RECT  8.030 1.745 9.305 1.975 ;
        RECT  8.070 2.895 9.305 3.125 ;
        RECT  7.840 2.895 8.070 3.835 ;
        RECT  7.800 1.370 8.030 1.975 ;
        RECT  7.570 0.740 7.930 0.970 ;
        RECT  7.730 3.460 7.840 3.835 ;
        RECT  6.550 3.605 7.730 3.835 ;
        RECT  7.340 0.740 7.570 1.365 ;
        RECT  7.295 2.460 7.390 2.800 ;
        RECT  7.295 1.635 7.350 1.975 ;
        RECT  5.665 1.135 7.340 1.365 ;
        RECT  7.065 1.635 7.295 3.375 ;
        RECT  7.010 1.635 7.065 1.975 ;
        RECT  7.010 2.460 7.065 3.375 ;
        RECT  6.780 2.905 7.010 3.375 ;
        RECT  6.095 2.905 6.780 3.135 ;
        RECT  6.320 3.545 6.550 3.835 ;
        RECT  3.715 3.545 6.320 3.775 ;
        RECT  5.865 2.540 6.095 3.135 ;
        RECT  5.635 1.120 5.665 1.460 ;
        RECT  5.405 1.120 5.635 3.135 ;
        RECT  5.325 1.120 5.405 1.460 ;
        RECT  5.085 2.905 5.405 3.135 ;
        RECT  4.930 1.840 5.160 2.205 ;
        RECT  4.040 2.905 5.085 3.260 ;
        RECT  3.580 1.975 4.930 2.205 ;
        RECT  3.810 2.510 4.040 3.260 ;
        RECT  3.485 3.545 3.715 4.365 ;
        RECT  3.350 0.955 3.580 2.965 ;
        RECT  3.135 4.135 3.485 4.365 ;
        RECT  3.025 0.955 3.350 1.240 ;
        RECT  3.050 2.735 3.350 2.965 ;
        RECT  2.890 1.770 3.120 2.225 ;
        RECT  2.820 2.735 3.050 3.820 ;
        RECT  2.685 0.900 3.025 1.240 ;
        RECT  2.425 1.995 2.890 2.225 ;
        RECT  2.425 3.280 2.500 3.645 ;
        RECT  2.225 1.455 2.425 3.645 ;
        RECT  2.210 1.400 2.225 3.645 ;
        RECT  1.870 0.640 2.220 1.050 ;
        RECT  2.195 1.400 2.210 3.535 ;
        RECT  1.885 1.400 2.195 1.740 ;
        RECT  1.550 3.250 2.195 3.535 ;
        RECT  1.735 3.970 2.075 4.310 ;
        RECT  0.520 0.820 1.870 1.050 ;
        RECT  0.465 3.980 1.735 4.210 ;
        RECT  0.290 0.820 0.520 1.745 ;
        RECT  0.465 3.270 0.520 3.610 ;
        RECT  0.235 3.270 0.465 4.210 ;
        RECT  0.180 1.405 0.290 1.745 ;
        RECT  0.180 3.270 0.235 3.610 ;
    END
END DFFSRX1

MACRO DFFSHQXL
    CLASS CORE ;
    FOREIGN DFFSHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.005 2.190 11.305 2.530 ;
        RECT  10.965 2.190 11.005 2.635 ;
        RECT  10.855 2.220 10.965 2.635 ;
        RECT  10.625 2.220 10.855 4.175 ;
        RECT  5.415 3.945 10.625 4.175 ;
        RECT  5.185 2.660 5.415 4.175 ;
        RECT  5.065 2.660 5.185 2.945 ;
        RECT  4.835 2.405 5.065 2.945 ;
        RECT  4.165 2.555 4.835 2.945 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 1.120 12.985 3.005 ;
        RECT  12.495 1.120 12.755 1.460 ;
        RECT  12.680 2.635 12.755 3.005 ;
        RECT  11.825 2.775 12.680 3.005 ;
        RECT  11.595 2.775 11.825 3.460 ;
        RECT  11.485 3.120 11.595 3.460 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.855 1.840 2.480 ;
        RECT  1.365 1.805 1.765 2.480 ;
        RECT  1.280 1.855 1.365 2.480 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 0.635 0.770 1.095 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.555 -0.400 13.200 0.400 ;
        RECT  11.215 -0.400 11.555 1.430 ;
        RECT  9.850 -0.400 11.215 0.400 ;
        RECT  9.510 -0.400 9.850 0.575 ;
        RECT  6.865 -0.400 9.510 0.400 ;
        RECT  6.635 -0.400 6.865 1.495 ;
        RECT  4.040 -0.400 6.635 0.400 ;
        RECT  3.700 -0.400 4.040 0.845 ;
        RECT  1.355 -0.400 3.700 0.400 ;
        RECT  1.015 -0.400 1.355 0.575 ;
        RECT  0.000 -0.400 1.015 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.545 4.640 13.200 5.440 ;
        RECT  12.205 3.320 12.545 5.440 ;
        RECT  11.215 4.640 12.205 5.440 ;
        RECT  10.875 4.465 11.215 5.440 ;
        RECT  9.835 4.640 10.875 5.440 ;
        RECT  9.495 4.465 9.835 5.440 ;
        RECT  6.660 4.640 9.495 5.440 ;
        RECT  6.295 4.465 6.660 5.440 ;
        RECT  4.950 4.640 6.295 5.440 ;
        RECT  4.010 4.140 4.950 5.440 ;
        RECT  1.450 4.640 4.010 5.440 ;
        RECT  1.110 4.465 1.450 5.440 ;
        RECT  0.000 4.640 1.110 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.440 2.165 12.445 2.450 ;
        RECT  12.215 1.725 12.440 2.450 ;
        RECT  12.210 1.725 12.215 2.395 ;
        RECT  10.605 1.725 12.210 1.955 ;
        RECT  10.490 0.805 10.605 1.955 ;
        RECT  10.375 0.695 10.490 1.955 ;
        RECT  10.135 0.695 10.375 1.040 ;
        RECT  10.140 2.640 10.345 3.150 ;
        RECT  10.115 1.290 10.140 3.150 ;
        RECT  9.560 0.810 10.135 1.040 ;
        RECT  9.910 1.290 10.115 2.870 ;
        RECT  9.250 2.640 9.910 2.870 ;
        RECT  9.330 0.810 9.560 2.265 ;
        RECT  8.485 0.810 9.330 1.040 ;
        RECT  8.790 2.035 9.330 2.265 ;
        RECT  9.020 2.640 9.250 3.000 ;
        RECT  8.330 1.485 8.900 1.715 ;
        RECT  6.725 3.440 8.865 3.670 ;
        RECT  8.560 2.035 8.790 3.190 ;
        RECT  7.920 2.960 8.560 3.190 ;
        RECT  8.145 0.755 8.485 1.095 ;
        RECT  8.100 1.485 8.330 2.445 ;
        RECT  7.710 2.215 8.100 2.445 ;
        RECT  7.615 1.105 7.725 1.445 ;
        RECT  7.480 2.215 7.710 2.580 ;
        RECT  7.385 1.105 7.615 1.965 ;
        RECT  7.235 2.960 7.410 3.190 ;
        RECT  7.235 1.735 7.385 1.965 ;
        RECT  7.005 1.735 7.235 3.190 ;
        RECT  6.495 1.870 6.725 3.670 ;
        RECT  6.395 1.870 6.495 2.100 ;
        RECT  6.375 3.395 6.495 3.670 ;
        RECT  6.165 1.350 6.395 2.100 ;
        RECT  5.645 3.395 6.375 3.625 ;
        RECT  5.935 2.330 6.260 2.670 ;
        RECT  6.065 1.350 6.165 1.580 ;
        RECT  5.835 0.675 6.065 1.580 ;
        RECT  5.920 1.810 5.935 2.670 ;
        RECT  5.705 1.810 5.920 2.615 ;
        RECT  5.500 0.675 5.835 0.905 ;
        RECT  5.550 1.810 5.705 2.040 ;
        RECT  5.320 1.335 5.550 2.040 ;
        RECT  4.960 1.335 5.320 1.995 ;
        RECT  4.625 0.775 5.065 1.005 ;
        RECT  3.935 1.765 4.960 1.995 ;
        RECT  4.320 3.340 4.660 3.680 ;
        RECT  4.395 0.775 4.625 1.365 ;
        RECT  2.990 1.135 4.395 1.365 ;
        RECT  3.935 3.340 4.320 3.570 ;
        RECT  3.705 1.765 3.935 3.570 ;
        RECT  3.315 1.885 3.705 2.115 ;
        RECT  3.245 2.360 3.475 3.635 ;
        RECT  2.985 2.360 3.245 2.590 ;
        RECT  2.775 3.405 3.245 3.635 ;
        RECT  2.340 2.870 3.015 3.100 ;
        RECT  2.985 1.015 2.990 1.365 ;
        RECT  2.755 1.015 2.985 2.590 ;
        RECT  2.435 3.405 2.775 3.745 ;
        RECT  2.675 1.015 2.755 1.300 ;
        RECT  2.335 0.960 2.675 1.300 ;
        RECT  2.110 1.715 2.340 3.100 ;
        RECT  0.890 2.870 2.110 3.100 ;
        RECT  0.590 2.870 0.890 3.490 ;
        RECT  0.590 1.345 0.645 1.685 ;
        RECT  0.550 1.345 0.590 3.490 ;
        RECT  0.360 1.345 0.550 3.100 ;
        RECT  0.305 1.345 0.360 1.685 ;
    END
END DFFSHQXL

MACRO DFFSHQX4
    CLASS CORE ;
    FOREIGN DFFSHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSHQXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.715 2.250 16.940 2.480 ;
        RECT  16.380 2.250 16.715 2.565 ;
        RECT  15.055 2.335 16.380 2.565 ;
        RECT  15.010 2.255 15.055 2.565 ;
        RECT  14.780 2.255 15.010 4.235 ;
        RECT  14.640 2.255 14.780 2.485 ;
        RECT  14.660 3.755 14.780 4.235 ;
        RECT  10.045 4.005 14.660 4.235 ;
        RECT  9.815 3.530 10.045 4.235 ;
        RECT  5.645 3.530 9.815 3.760 ;
        RECT  5.645 2.965 5.725 3.195 ;
        RECT  5.415 2.900 5.645 3.760 ;
        RECT  4.430 2.900 5.415 3.130 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.280 0.800 18.300 1.290 ;
        RECT  18.050 0.800 18.280 3.185 ;
        RECT  17.960 0.800 18.050 1.495 ;
        RECT  17.680 2.955 18.050 3.185 ;
        RECT  15.740 1.265 17.960 1.495 ;
        RECT  17.300 2.940 17.680 4.340 ;
        RECT  17.080 2.985 17.300 4.030 ;
        RECT  17.020 2.985 17.080 3.220 ;
        RECT  15.980 2.985 17.020 3.215 ;
        RECT  15.900 2.985 15.980 3.220 ;
        RECT  15.560 2.985 15.900 3.925 ;
        RECT  15.505 1.055 15.740 1.495 ;
        RECT  15.400 1.055 15.505 1.395 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.375 1.955 2.875 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.820 1.180 2.545 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.020 -0.400 18.480 0.400 ;
        RECT  16.680 -0.400 17.020 0.955 ;
        RECT  14.250 -0.400 16.680 0.400 ;
        RECT  12.970 -0.400 14.250 0.575 ;
        RECT  8.820 -0.400 12.970 0.400 ;
        RECT  8.480 -0.400 8.820 1.280 ;
        RECT  7.375 -0.400 8.480 0.400 ;
        RECT  7.035 -0.400 7.375 1.395 ;
        RECT  4.085 -0.400 7.035 0.400 ;
        RECT  3.745 -0.400 4.085 0.575 ;
        RECT  1.520 -0.400 3.745 0.400 ;
        RECT  1.180 -0.400 1.520 0.575 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.215 4.640 18.480 5.440 ;
        RECT  17.985 3.480 18.215 5.440 ;
        RECT  16.660 4.640 17.985 5.440 ;
        RECT  16.320 3.480 16.660 5.440 ;
        RECT  15.100 4.640 16.320 5.440 ;
        RECT  14.760 4.465 15.100 5.440 ;
        RECT  13.630 4.640 14.760 5.440 ;
        RECT  13.290 4.465 13.630 5.440 ;
        RECT  8.950 4.640 13.290 5.440 ;
        RECT  8.610 4.465 8.950 5.440 ;
        RECT  7.425 4.640 8.610 5.440 ;
        RECT  7.085 4.465 7.425 5.440 ;
        RECT  5.960 4.640 7.085 5.440 ;
        RECT  5.620 4.465 5.960 5.440 ;
        RECT  4.440 4.640 5.620 5.440 ;
        RECT  4.100 4.465 4.440 5.440 ;
        RECT  1.730 4.640 4.100 5.440 ;
        RECT  1.390 4.465 1.730 5.440 ;
        RECT  0.000 4.640 1.390 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.710 2.205 17.820 2.545 ;
        RECT  17.480 1.780 17.710 2.545 ;
        RECT  16.080 1.780 17.480 2.010 ;
        RECT  15.680 1.780 16.080 2.065 ;
        RECT  15.015 1.780 15.680 2.010 ;
        RECT  14.785 0.865 15.015 2.010 ;
        RECT  12.205 0.865 14.785 1.095 ;
        RECT  14.310 3.000 14.420 3.340 ;
        RECT  14.080 1.545 14.310 3.340 ;
        RECT  13.260 1.545 14.080 1.775 ;
        RECT  13.705 2.250 13.815 2.590 ;
        RECT  13.475 2.250 13.705 3.775 ;
        RECT  12.205 3.545 13.475 3.775 ;
        RECT  12.920 1.370 13.260 1.775 ;
        RECT  12.885 1.540 12.920 1.775 ;
        RECT  12.600 1.540 12.885 2.345 ;
        RECT  12.545 2.005 12.600 2.345 ;
        RECT  11.975 0.865 12.205 3.775 ;
        RECT  11.700 0.865 11.975 1.095 ;
        RECT  10.420 3.545 11.975 3.775 ;
        RECT  11.590 0.865 11.700 1.410 ;
        RECT  11.360 0.725 11.590 1.410 ;
        RECT  10.880 3.070 11.520 3.300 ;
        RECT  10.260 0.725 11.360 0.955 ;
        RECT  10.880 1.200 10.980 1.540 ;
        RECT  10.650 1.200 10.880 3.300 ;
        RECT  10.640 1.200 10.650 1.745 ;
        RECT  7.845 3.070 10.650 3.300 ;
        RECT  9.540 1.515 10.640 1.745 ;
        RECT  10.030 0.725 10.260 1.280 ;
        RECT  9.920 0.940 10.030 1.280 ;
        RECT  7.585 1.975 10.025 2.205 ;
        RECT  9.200 1.100 9.540 1.745 ;
        RECT  9.255 3.995 9.485 4.405 ;
        RECT  3.495 3.995 9.255 4.225 ;
        RECT  8.100 1.515 9.200 1.745 ;
        RECT  7.815 1.110 8.100 1.745 ;
        RECT  7.760 1.110 7.815 1.450 ;
        RECT  7.355 1.725 7.585 3.155 ;
        RECT  6.585 1.725 7.355 1.955 ;
        RECT  6.465 2.925 7.355 3.155 ;
        RECT  5.635 2.260 7.120 2.490 ;
        RECT  6.355 0.775 6.585 1.955 ;
        RECT  4.850 0.775 6.355 1.005 ;
        RECT  5.565 1.300 5.635 2.665 ;
        RECT  5.405 1.245 5.565 2.665 ;
        RECT  5.225 1.245 5.405 1.585 ;
        RECT  3.865 2.435 5.405 2.665 ;
        RECT  3.200 1.975 5.175 2.205 ;
        RECT  4.915 3.365 5.145 3.760 ;
        RECT  3.865 3.365 4.915 3.595 ;
        RECT  4.620 0.775 4.850 1.705 ;
        RECT  3.485 1.475 4.620 1.705 ;
        RECT  3.635 2.435 3.865 3.595 ;
        RECT  3.210 3.995 3.495 4.235 ;
        RECT  3.255 0.635 3.485 1.705 ;
        RECT  3.075 0.635 3.255 0.865 ;
        RECT  2.735 4.005 3.210 4.235 ;
        RECT  3.020 1.975 3.200 3.715 ;
        RECT  2.970 1.175 3.020 3.715 ;
        RECT  2.790 1.175 2.970 2.205 ;
        RECT  2.500 1.175 2.790 1.405 ;
        RECT  2.505 3.605 2.735 4.235 ;
        RECT  2.415 3.605 2.505 3.835 ;
        RECT  2.185 1.740 2.415 3.835 ;
        RECT  0.955 3.605 2.185 3.835 ;
        RECT  0.615 3.000 0.955 3.940 ;
        RECT  0.570 1.180 0.760 1.520 ;
        RECT  0.570 3.000 0.615 3.230 ;
        RECT  0.420 1.180 0.570 3.230 ;
        RECT  0.340 1.235 0.420 3.230 ;
    END
END DFFSHQX4

MACRO DFFSHQX2
    CLASS CORE ;
    FOREIGN DFFSHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSHQXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.160 2.110 15.215 2.450 ;
        RECT  14.930 2.110 15.160 3.755 ;
        RECT  14.875 2.110 14.930 2.450 ;
        RECT  12.755 3.525 14.930 3.755 ;
        RECT  12.550 2.175 12.780 2.515 ;
        RECT  12.550 3.500 12.755 3.755 ;
        RECT  12.440 2.175 12.550 3.755 ;
        RECT  12.410 2.230 12.440 3.755 ;
        RECT  12.320 2.230 12.410 4.305 ;
        RECT  12.180 3.525 12.320 4.305 ;
        RECT  8.360 4.075 12.180 4.305 ;
        RECT  8.130 3.655 8.360 4.305 ;
        RECT  8.060 3.655 8.130 4.085 ;
        RECT  7.120 3.655 8.060 3.885 ;
        RECT  6.930 3.655 7.120 4.085 ;
        RECT  6.700 3.655 6.930 4.365 ;
        RECT  5.145 4.135 6.700 4.365 ;
        RECT  5.065 2.455 5.145 4.365 ;
        RECT  4.915 2.405 5.065 4.365 ;
        RECT  4.115 2.405 4.915 2.685 ;
        RECT  3.830 2.405 4.115 2.780 ;
        RECT  3.775 2.440 3.830 2.780 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.415 1.315 14.645 3.080 ;
        RECT  14.210 1.315 14.415 1.545 ;
        RECT  14.075 2.850 14.415 3.080 ;
        RECT  13.870 1.205 14.210 1.545 ;
        RECT  13.740 2.850 14.075 3.190 ;
        RECT  13.415 2.850 13.740 3.195 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.055 1.820 1.475 2.755 ;
        RECT  0.875 1.845 1.055 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 3.805 0.675 4.235 ;
        RECT  0.215 3.805 0.475 4.315 ;
        RECT  0.190 3.805 0.215 4.235 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.490 -0.400 15.840 0.400 ;
        RECT  15.150 -0.400 15.490 1.510 ;
        RECT  12.410 -0.400 15.150 0.400 ;
        RECT  12.070 -0.400 12.410 0.575 ;
        RECT  8.285 -0.400 12.070 0.400 ;
        RECT  7.945 -0.400 8.285 1.390 ;
        RECT  6.790 -0.400 7.945 0.400 ;
        RECT  6.560 -0.400 6.790 1.370 ;
        RECT  3.865 -0.400 6.560 0.400 ;
        RECT  3.525 -0.400 3.865 0.960 ;
        RECT  1.280 -0.400 3.525 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.515 4.640 15.840 5.440 ;
        RECT  14.175 4.085 14.515 5.440 ;
        RECT  13.015 4.640 14.175 5.440 ;
        RECT  12.675 4.035 13.015 5.440 ;
        RECT  7.750 4.640 12.675 5.440 ;
        RECT  7.410 4.170 7.750 5.440 ;
        RECT  4.545 4.640 7.410 5.440 ;
        RECT  3.735 4.140 4.545 5.440 ;
        RECT  1.310 4.640 3.735 5.440 ;
        RECT  0.970 4.465 1.310 5.440 ;
        RECT  0.000 4.640 0.970 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.725 2.040 14.065 2.380 ;
        RECT  13.250 2.040 13.725 2.270 ;
        RECT  13.020 0.865 13.250 2.270 ;
        RECT  10.475 0.865 13.020 1.095 ;
        RECT  11.720 2.125 11.950 3.745 ;
        RECT  11.645 2.125 11.720 2.355 ;
        RECT  11.430 3.515 11.720 3.745 ;
        RECT  11.645 1.460 11.700 1.800 ;
        RECT  11.415 1.460 11.645 2.355 ;
        RECT  10.475 2.815 11.485 3.045 ;
        RECT  11.360 1.460 11.415 1.800 ;
        RECT  11.400 2.060 11.415 2.355 ;
        RECT  11.060 2.060 11.400 2.400 ;
        RECT  10.315 0.865 10.475 3.845 ;
        RECT  10.245 0.795 10.315 3.845 ;
        RECT  10.085 0.795 10.245 1.600 ;
        RECT  8.890 3.615 10.245 3.845 ;
        RECT  8.985 0.795 10.085 1.025 ;
        RECT  9.755 3.135 10.010 3.365 ;
        RECT  9.705 1.625 9.755 3.365 ;
        RECT  9.525 1.280 9.705 3.365 ;
        RECT  9.365 1.280 9.525 1.860 ;
        RECT  6.695 3.135 9.525 3.365 ;
        RECT  7.565 1.630 9.365 1.860 ;
        RECT  6.465 2.090 9.285 2.320 ;
        RECT  8.755 0.795 8.985 1.280 ;
        RECT  8.645 0.940 8.755 1.280 ;
        RECT  7.335 1.115 7.565 1.860 ;
        RECT  7.225 1.115 7.335 1.455 ;
        RECT  6.235 1.750 6.465 3.845 ;
        RECT  6.090 1.750 6.235 1.980 ;
        RECT  5.845 3.560 6.235 3.845 ;
        RECT  5.990 1.410 6.090 1.980 ;
        RECT  5.860 0.675 5.990 1.980 ;
        RECT  5.750 2.240 5.980 2.875 ;
        RECT  5.760 0.675 5.860 1.640 ;
        RECT  5.505 3.560 5.845 3.900 ;
        RECT  5.345 0.675 5.760 0.905 ;
        RECT  5.620 2.240 5.750 2.470 ;
        RECT  5.390 1.875 5.620 2.470 ;
        RECT  5.245 1.875 5.390 2.105 ;
        RECT  5.015 1.415 5.245 2.105 ;
        RECT  4.905 1.415 5.015 1.885 ;
        RECT  4.665 0.720 5.005 1.060 ;
        RECT  3.440 1.655 4.905 1.885 ;
        RECT  4.545 0.830 4.665 1.060 ;
        RECT  4.315 0.830 4.545 1.420 ;
        RECT  4.180 3.300 4.520 3.640 ;
        RECT  2.620 1.190 4.315 1.420 ;
        RECT  3.385 3.355 4.180 3.585 ;
        RECT  3.385 1.655 3.440 2.510 ;
        RECT  3.210 1.655 3.385 3.585 ;
        RECT  3.155 2.170 3.210 3.585 ;
        RECT  3.100 2.170 3.155 2.510 ;
        RECT  2.120 3.960 2.975 4.190 ;
        RECT  2.390 1.190 2.620 3.570 ;
        RECT  2.350 1.190 2.390 1.585 ;
        RECT  2.350 3.135 2.390 3.570 ;
        RECT  2.140 1.355 2.350 1.585 ;
        RECT  2.120 1.835 2.155 2.205 ;
        RECT  1.890 1.835 2.120 4.190 ;
        RECT  0.615 3.245 1.890 3.475 ;
        RECT  0.375 3.135 0.615 3.475 ;
        RECT  0.375 1.455 0.560 1.795 ;
        RECT  0.145 1.455 0.375 3.475 ;
    END
END DFFSHQX2

MACRO DFFSHQX1
    CLASS CORE ;
    FOREIGN DFFSHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSHQXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.435 1.845 11.665 2.100 ;
        RECT  11.305 1.870 11.435 2.100 ;
        RECT  11.075 1.870 11.305 2.450 ;
        RECT  10.965 2.110 11.075 2.450 ;
        RECT  10.855 2.220 10.965 2.450 ;
        RECT  10.625 2.220 10.855 4.175 ;
        RECT  5.415 3.945 10.625 4.175 ;
        RECT  5.185 2.660 5.415 4.175 ;
        RECT  5.065 2.660 5.185 2.945 ;
        RECT  4.835 2.405 5.065 2.945 ;
        RECT  4.165 2.555 4.835 2.945 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 0.855 12.985 3.005 ;
        RECT  12.680 0.855 12.755 1.285 ;
        RECT  12.680 2.635 12.755 3.005 ;
        RECT  12.550 0.855 12.680 1.220 ;
        RECT  11.825 2.775 12.680 3.005 ;
        RECT  11.595 2.775 11.825 3.440 ;
        RECT  11.485 3.100 11.595 3.440 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 1.820 1.840 2.380 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.675 1.180 3.220 ;
        RECT  0.605 2.675 0.800 3.055 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.595 -0.400 13.200 0.400 ;
        RECT  11.175 -0.400 11.595 1.010 ;
        RECT  9.850 -0.400 11.175 0.400 ;
        RECT  9.510 -0.400 9.850 0.575 ;
        RECT  6.865 -0.400 9.510 0.400 ;
        RECT  6.635 -0.400 6.865 1.280 ;
        RECT  4.040 -0.400 6.635 0.400 ;
        RECT  3.700 -0.400 4.040 0.845 ;
        RECT  1.280 -0.400 3.700 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.545 4.640 13.200 5.440 ;
        RECT  12.205 3.320 12.545 5.440 ;
        RECT  11.240 4.640 12.205 5.440 ;
        RECT  10.900 4.465 11.240 5.440 ;
        RECT  9.835 4.640 10.900 5.440 ;
        RECT  9.495 4.465 9.835 5.440 ;
        RECT  6.660 4.640 9.495 5.440 ;
        RECT  6.295 4.465 6.660 5.440 ;
        RECT  4.950 4.640 6.295 5.440 ;
        RECT  4.010 4.140 4.950 5.440 ;
        RECT  1.100 4.640 4.010 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.260 2.165 12.420 2.395 ;
        RECT  12.030 1.285 12.260 2.395 ;
        RECT  10.605 1.285 12.030 1.515 ;
        RECT  10.490 0.805 10.605 1.515 ;
        RECT  10.375 0.695 10.490 1.515 ;
        RECT  10.155 2.640 10.385 3.150 ;
        RECT  10.135 0.695 10.375 1.035 ;
        RECT  10.140 2.640 10.155 2.870 ;
        RECT  9.910 1.320 10.140 2.870 ;
        RECT  9.380 0.805 10.135 1.035 ;
        RECT  9.250 2.640 9.910 2.870 ;
        RECT  9.150 0.805 9.380 2.265 ;
        RECT  9.020 2.640 9.250 3.000 ;
        RECT  8.665 0.805 9.150 1.035 ;
        RECT  8.790 2.035 9.150 2.265 ;
        RECT  8.330 1.450 8.900 1.680 ;
        RECT  6.725 3.440 8.865 3.670 ;
        RECT  8.560 2.035 8.790 3.190 ;
        RECT  8.430 0.805 8.665 1.220 ;
        RECT  7.920 2.960 8.560 3.190 ;
        RECT  8.025 0.990 8.430 1.220 ;
        RECT  8.100 1.450 8.330 2.445 ;
        RECT  7.710 2.215 8.100 2.445 ;
        RECT  7.480 2.215 7.710 2.580 ;
        RECT  7.530 1.080 7.640 1.420 ;
        RECT  7.300 1.080 7.530 1.835 ;
        RECT  7.235 2.960 7.455 3.190 ;
        RECT  7.235 1.605 7.300 1.835 ;
        RECT  7.005 1.605 7.235 3.190 ;
        RECT  6.495 1.595 6.725 3.670 ;
        RECT  6.395 1.595 6.495 1.825 ;
        RECT  6.375 3.385 6.495 3.670 ;
        RECT  6.165 1.350 6.395 1.825 ;
        RECT  5.685 3.385 6.375 3.615 ;
        RECT  5.935 2.355 6.260 2.585 ;
        RECT  6.065 1.350 6.165 1.580 ;
        RECT  5.835 0.675 6.065 1.580 ;
        RECT  5.705 1.810 5.935 2.585 ;
        RECT  5.500 0.675 5.835 0.905 ;
        RECT  5.550 1.810 5.705 2.040 ;
        RECT  5.320 1.335 5.550 2.040 ;
        RECT  4.960 1.335 5.320 1.995 ;
        RECT  4.625 0.775 5.065 1.005 ;
        RECT  3.935 1.765 4.960 1.995 ;
        RECT  3.935 3.395 4.660 3.625 ;
        RECT  4.395 0.775 4.625 1.365 ;
        RECT  2.990 1.135 4.395 1.365 ;
        RECT  3.705 1.765 3.935 3.625 ;
        RECT  3.315 1.845 3.705 2.075 ;
        RECT  3.245 2.365 3.475 3.890 ;
        RECT  2.985 2.365 3.245 2.595 ;
        RECT  2.385 3.660 3.245 3.890 ;
        RECT  2.985 0.855 2.990 1.365 ;
        RECT  2.755 0.855 2.985 2.595 ;
        RECT  2.345 2.995 2.965 3.225 ;
        RECT  2.335 0.855 2.755 1.085 ;
        RECT  2.115 1.775 2.345 3.425 ;
        RECT  1.820 3.195 2.115 3.425 ;
        RECT  1.590 3.195 1.820 3.870 ;
        RECT  0.520 3.640 1.590 3.870 ;
        RECT  0.370 3.320 0.520 3.870 ;
        RECT  0.370 1.385 0.465 1.755 ;
        RECT  0.140 1.385 0.370 3.870 ;
    END
END DFFSHQX1

MACRO DFFSXL
    CLASS CORE ;
    FOREIGN DFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 3.900 9.790 4.410 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.460 0.870 11.690 3.970 ;
        RECT  10.945 0.870 11.460 1.100 ;
        RECT  11.100 3.740 11.460 3.970 ;
        RECT  11.005 3.740 11.100 4.210 ;
        RECT  10.760 3.740 11.005 4.315 ;
        RECT  10.605 0.755 10.945 1.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.325 3.090 12.360 3.430 ;
        RECT  12.095 1.250 12.325 3.430 ;
        RECT  11.960 1.250 12.095 1.590 ;
        RECT  12.020 3.090 12.095 3.430 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 1.205 1.835 1.705 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.030 2.965 1.105 3.195 ;
        RECT  0.800 2.480 1.030 3.195 ;
        RECT  0.605 2.480 0.800 2.820 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.165 -0.400 12.540 0.400 ;
        RECT  11.825 -0.400 12.165 0.575 ;
        RECT  10.220 -0.400 11.825 0.400 ;
        RECT  9.880 -0.400 10.220 1.095 ;
        RECT  8.560 -0.400 9.880 0.400 ;
        RECT  8.220 -0.400 8.560 0.575 ;
        RECT  6.165 -0.400 8.220 0.400 ;
        RECT  5.935 -0.400 6.165 1.010 ;
        RECT  4.040 -0.400 5.935 0.400 ;
        RECT  3.700 -0.400 4.040 1.090 ;
        RECT  1.535 -0.400 3.700 0.400 ;
        RECT  1.195 -0.400 1.535 0.575 ;
        RECT  0.000 -0.400 1.195 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 4.640 12.540 5.440 ;
        RECT  12.305 4.465 12.360 5.440 ;
        RECT  12.075 4.410 12.305 5.440 ;
        RECT  12.020 4.465 12.075 5.440 ;
        RECT  10.380 4.640 12.020 5.440 ;
        RECT  10.040 3.170 10.380 5.440 ;
        RECT  8.930 4.640 10.040 5.440 ;
        RECT  8.590 4.080 8.930 5.440 ;
        RECT  6.420 4.640 8.590 5.440 ;
        RECT  6.080 4.135 6.420 5.440 ;
        RECT  5.160 4.640 6.080 5.440 ;
        RECT  4.820 4.135 5.160 5.440 ;
        RECT  3.760 4.640 4.820 5.440 ;
        RECT  3.420 4.465 3.760 5.440 ;
        RECT  1.300 4.640 3.420 5.440 ;
        RECT  0.960 4.465 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.100 2.110 11.225 2.450 ;
        RECT  10.985 1.570 11.100 3.510 ;
        RECT  10.870 1.460 10.985 3.510 ;
        RECT  10.645 1.460 10.870 1.800 ;
        RECT  10.760 3.170 10.870 3.510 ;
        RECT  9.660 1.985 10.370 2.325 ;
        RECT  9.430 1.455 9.660 3.510 ;
        RECT  7.880 1.455 9.430 1.685 ;
        RECT  9.320 3.170 9.430 3.510 ;
        RECT  8.390 2.410 9.200 2.750 ;
        RECT  8.160 1.915 8.390 3.210 ;
        RECT  7.325 1.915 8.160 2.145 ;
        RECT  7.740 2.980 8.160 3.210 ;
        RECT  6.840 2.500 7.930 2.730 ;
        RECT  7.400 2.980 7.740 3.320 ;
        RECT  7.260 3.930 7.370 4.270 ;
        RECT  7.095 1.470 7.325 2.145 ;
        RECT  7.030 3.675 7.260 4.270 ;
        RECT  5.730 3.675 7.030 3.905 ;
        RECT  6.610 1.240 6.840 3.330 ;
        RECT  5.705 1.240 6.610 1.470 ;
        RECT  5.920 3.100 6.610 3.330 ;
        RECT  5.245 2.165 6.375 2.505 ;
        RECT  5.580 3.100 5.920 3.440 ;
        RECT  5.390 3.675 5.730 3.945 ;
        RECT  5.475 0.780 5.705 1.470 ;
        RECT  5.385 0.780 5.475 1.010 ;
        RECT  2.880 3.675 5.390 3.905 ;
        RECT  5.040 0.630 5.385 1.010 ;
        RECT  5.015 1.460 5.245 3.235 ;
        RECT  4.270 0.630 5.040 0.860 ;
        RECT  4.560 3.005 5.015 3.235 ;
        RECT  4.620 2.430 4.730 2.770 ;
        RECT  4.390 2.180 4.620 2.770 ;
        RECT  4.220 3.005 4.560 3.440 ;
        RECT  2.910 2.180 4.390 2.410 ;
        RECT  3.600 3.005 4.220 3.235 ;
        RECT  3.370 2.640 3.600 3.235 ;
        RECT  3.260 2.640 3.370 2.980 ;
        RECT  2.900 0.760 2.910 2.410 ;
        RECT  2.670 0.750 2.900 3.240 ;
        RECT  2.540 3.675 2.880 4.140 ;
        RECT  2.515 0.750 2.670 1.090 ;
        RECT  2.600 3.010 2.670 3.240 ;
        RECT  2.260 3.010 2.600 3.350 ;
        RECT  1.905 3.675 2.540 3.905 ;
        RECT  2.095 1.850 2.435 2.190 ;
        RECT  1.905 1.960 2.095 2.190 ;
        RECT  1.655 1.960 1.905 3.905 ;
        RECT  0.530 1.960 1.655 2.190 ;
        RECT  0.540 3.450 1.655 3.680 ;
        RECT  0.200 3.220 0.540 3.680 ;
        RECT  0.300 1.190 0.530 2.190 ;
        RECT  0.190 1.190 0.300 1.530 ;
    END
END DFFSXL

MACRO DFFSX4
    CLASS CORE ;
    FOREIGN DFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.260 4.050 5.140 4.410 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.210 1.820 16.360 3.220 ;
        RECT  16.060 1.260 16.210 3.220 ;
        RECT  15.980 0.855 16.060 3.220 ;
        RECT  15.720 0.855 15.980 1.665 ;
        RECT  15.600 2.780 15.980 3.120 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.960 1.820 18.340 3.220 ;
        RECT  17.500 1.820 17.960 2.050 ;
        RECT  17.325 2.985 17.960 3.215 ;
        RECT  17.270 0.855 17.500 2.050 ;
        RECT  17.095 2.985 17.325 3.975 ;
        RECT  17.160 0.855 17.270 1.665 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.820 1.845 2.100 ;
        RECT  1.305 1.670 1.840 2.140 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 2.380 1.180 2.660 ;
        RECT  0.605 2.210 0.945 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.220 -0.400 18.480 0.400 ;
        RECT  17.880 -0.400 18.220 1.485 ;
        RECT  16.780 -0.400 17.880 0.400 ;
        RECT  16.440 -0.400 16.780 1.485 ;
        RECT  15.340 -0.400 16.440 0.400 ;
        RECT  15.000 -0.400 15.340 0.950 ;
        RECT  14.040 -0.400 15.000 0.400 ;
        RECT  13.700 -0.400 14.040 1.550 ;
        RECT  11.440 -0.400 13.700 0.400 ;
        RECT  11.100 -0.400 11.440 0.575 ;
        RECT  9.450 -0.400 11.100 0.400 ;
        RECT  9.110 -0.400 9.450 1.320 ;
        RECT  6.890 -0.400 9.110 0.400 ;
        RECT  6.550 -0.400 6.890 1.320 ;
        RECT  3.970 -0.400 6.550 0.400 ;
        RECT  3.630 -0.400 3.970 1.280 ;
        RECT  1.250 -0.400 3.630 0.400 ;
        RECT  0.910 -0.400 1.250 0.575 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.100 4.640 18.480 5.440 ;
        RECT  17.760 3.605 18.100 5.440 ;
        RECT  16.660 4.640 17.760 5.440 ;
        RECT  16.320 4.030 16.660 5.440 ;
        RECT  15.220 4.640 16.320 5.440 ;
        RECT  14.880 4.090 15.220 5.440 ;
        RECT  13.960 4.640 14.880 5.440 ;
        RECT  13.620 2.975 13.960 5.440 ;
        RECT  12.520 4.640 13.620 5.440 ;
        RECT  12.180 3.435 12.520 5.440 ;
        RECT  11.040 4.640 12.180 5.440 ;
        RECT  10.700 4.040 11.040 5.440 ;
        RECT  9.330 4.640 10.700 5.440 ;
        RECT  8.990 3.600 9.330 5.440 ;
        RECT  6.780 4.640 8.990 5.440 ;
        RECT  6.440 4.140 6.780 5.440 ;
        RECT  5.600 4.640 6.440 5.440 ;
        RECT  5.370 4.140 5.600 5.440 ;
        RECT  4.030 4.640 5.370 5.440 ;
        RECT  3.690 4.150 4.030 5.440 ;
        RECT  1.265 4.640 3.690 5.440 ;
        RECT  0.925 4.465 1.265 5.440 ;
        RECT  0.000 4.640 0.925 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.860 2.040 17.030 2.380 ;
        RECT  16.630 2.040 16.860 3.685 ;
        RECT  14.760 3.455 16.630 3.685 ;
        RECT  14.760 1.310 14.800 1.650 ;
        RECT  14.680 1.310 14.760 3.685 ;
        RECT  14.530 1.310 14.680 3.710 ;
        RECT  14.460 1.310 14.530 1.650 ;
        RECT  14.340 2.900 14.530 3.710 ;
        RECT  13.240 2.080 14.300 2.420 ;
        RECT  13.010 1.375 13.240 3.785 ;
        RECT  12.760 1.375 13.010 1.605 ;
        RECT  12.900 2.975 13.010 3.785 ;
        RECT  11.800 2.975 12.900 3.205 ;
        RECT  12.420 0.790 12.760 1.605 ;
        RECT  12.180 1.895 12.520 2.705 ;
        RECT  11.110 1.110 12.420 1.340 ;
        RECT  10.105 2.185 12.180 2.415 ;
        RECT  11.460 2.975 11.800 3.785 ;
        RECT  10.450 3.365 11.460 3.595 ;
        RECT  10.770 1.000 11.110 1.340 ;
        RECT  10.220 3.365 10.450 4.040 ;
        RECT  10.110 3.700 10.220 4.040 ;
        RECT  10.105 1.430 10.160 1.770 ;
        RECT  9.880 1.430 10.105 3.130 ;
        RECT  9.875 1.430 9.880 3.240 ;
        RECT  9.820 1.430 9.875 1.780 ;
        RECT  9.540 2.900 9.875 3.240 ;
        RECT  8.875 1.550 9.820 1.780 ;
        RECT  9.305 2.330 9.645 2.670 ;
        RECT  8.010 2.900 9.540 3.130 ;
        RECT  8.360 2.330 9.305 2.560 ;
        RECT  8.645 1.190 8.875 1.780 ;
        RECT  8.170 1.190 8.645 1.420 ;
        RECT  8.130 1.720 8.360 2.560 ;
        RECT  7.830 1.080 8.170 1.420 ;
        RECT  8.020 1.720 8.130 2.060 ;
        RECT  6.835 1.775 8.020 2.005 ;
        RECT  7.670 2.865 8.010 3.675 ;
        RECT  7.355 2.365 7.690 2.595 ;
        RECT  7.125 2.365 7.355 3.780 ;
        RECT  6.165 3.550 7.125 3.780 ;
        RECT  6.605 1.765 6.835 3.210 ;
        RECT  6.090 1.765 6.605 2.005 ;
        RECT  6.110 2.980 6.605 3.210 ;
        RECT  6.035 2.270 6.375 2.610 ;
        RECT  5.935 3.550 6.165 4.025 ;
        RECT  5.770 2.980 6.110 3.320 ;
        RECT  5.980 1.160 6.090 2.005 ;
        RECT  5.340 2.325 6.035 2.555 ;
        RECT  5.805 0.685 5.980 2.005 ;
        RECT  2.105 3.550 5.935 3.780 ;
        RECT  5.750 0.685 5.805 1.500 ;
        RECT  5.600 0.685 5.750 0.915 ;
        RECT  5.110 0.955 5.340 3.210 ;
        RECT  4.910 0.955 5.110 1.300 ;
        RECT  4.790 2.980 5.110 3.210 ;
        RECT  4.540 1.605 4.880 1.945 ;
        RECT  4.450 2.980 4.790 3.320 ;
        RECT  2.980 1.660 4.540 1.890 ;
        RECT  3.695 2.980 4.450 3.210 ;
        RECT  3.690 2.325 3.695 3.210 ;
        RECT  3.465 2.215 3.690 3.210 ;
        RECT  3.350 2.215 3.465 2.555 ;
        RECT  2.750 1.040 2.980 3.135 ;
        RECT  2.270 1.040 2.750 1.380 ;
        RECT  2.565 2.905 2.750 3.135 ;
        RECT  2.335 2.905 2.565 3.300 ;
        RECT  2.175 1.610 2.405 2.660 ;
        RECT  2.105 2.430 2.175 2.660 ;
        RECT  1.875 2.430 2.105 3.780 ;
        RECT  0.610 3.070 1.875 3.300 ;
        RECT  0.375 1.255 0.690 1.595 ;
        RECT  0.375 2.960 0.610 3.300 ;
        RECT  0.145 1.255 0.375 3.300 ;
    END
END DFFSX4

MACRO DFFSX2
    CLASS CORE ;
    FOREIGN DFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.085 4.005 9.685 4.355 ;
        RECT  3.930 4.005 9.085 4.235 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.860 1.260 12.325 1.540 ;
        RECT  11.630 0.630 11.860 2.940 ;
        RECT  11.370 0.630 11.630 0.970 ;
        RECT  11.580 2.635 11.630 2.940 ;
        RECT  11.360 2.635 11.580 3.050 ;
        RECT  11.240 2.710 11.360 3.050 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.415 1.325 13.645 3.115 ;
        RECT  13.340 1.260 13.415 3.115 ;
        RECT  13.230 1.260 13.340 1.555 ;
        RECT  13.020 2.885 13.340 3.115 ;
        RECT  12.890 0.745 13.230 1.555 ;
        RECT  12.680 2.885 13.020 4.165 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 2.360 1.805 2.755 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.135 2.295 0.515 2.830 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.470 -0.400 13.860 0.400 ;
        RECT  12.130 -0.400 12.470 0.575 ;
        RECT  11.010 -0.400 12.130 0.400 ;
        RECT  10.670 -0.400 11.010 0.575 ;
        RECT  8.630 -0.400 10.670 0.400 ;
        RECT  8.290 -0.400 8.630 1.565 ;
        RECT  6.085 -0.400 8.290 0.400 ;
        RECT  5.855 -0.400 6.085 1.300 ;
        RECT  3.860 -0.400 5.855 0.400 ;
        RECT  3.520 -0.400 3.860 1.130 ;
        RECT  1.450 -0.400 3.520 0.400 ;
        RECT  1.110 -0.400 1.450 0.575 ;
        RECT  0.000 -0.400 1.110 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.300 4.640 13.860 5.440 ;
        RECT  11.960 3.865 12.300 5.440 ;
        RECT  10.330 4.640 11.960 5.440 ;
        RECT  9.990 3.445 10.330 5.440 ;
        RECT  9.980 3.445 9.990 3.785 ;
        RECT  8.840 4.640 9.990 5.440 ;
        RECT  8.500 4.465 8.840 5.440 ;
        RECT  6.360 4.640 8.500 5.440 ;
        RECT  6.020 4.465 6.360 5.440 ;
        RECT  5.100 4.640 6.020 5.440 ;
        RECT  4.760 4.465 5.100 5.440 ;
        RECT  3.700 4.640 4.760 5.440 ;
        RECT  3.360 4.465 3.700 5.440 ;
        RECT  1.310 4.640 3.360 5.440 ;
        RECT  0.970 4.465 1.310 5.440 ;
        RECT  0.000 4.640 0.970 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.450 2.070 12.670 2.410 ;
        RECT  12.220 2.070 12.450 3.545 ;
        RECT  11.040 3.315 12.220 3.545 ;
        RECT  11.010 1.345 11.170 1.685 ;
        RECT  11.010 3.315 11.040 3.780 ;
        RECT  10.780 1.345 11.010 3.780 ;
        RECT  10.700 3.440 10.780 3.780 ;
        RECT  10.405 2.015 10.515 2.355 ;
        RECT  10.175 1.795 10.405 3.125 ;
        RECT  9.910 1.795 10.175 2.025 ;
        RECT  9.600 2.895 10.175 3.125 ;
        RECT  9.570 1.335 9.910 2.025 ;
        RECT  9.500 2.255 9.840 2.665 ;
        RECT  9.260 2.895 9.600 3.705 ;
        RECT  8.330 1.795 9.570 2.025 ;
        RECT  7.680 2.435 9.500 2.665 ;
        RECT  7.990 1.795 8.330 2.205 ;
        RECT  7.625 2.435 7.680 3.775 ;
        RECT  7.395 1.405 7.625 3.775 ;
        RECT  7.305 1.405 7.395 1.750 ;
        RECT  7.340 3.545 7.395 3.775 ;
        RECT  7.110 2.540 7.145 2.880 ;
        RECT  6.880 2.540 7.110 3.775 ;
        RECT  6.645 1.735 7.060 2.075 ;
        RECT  2.820 3.545 6.880 3.775 ;
        RECT  6.415 1.530 6.645 3.030 ;
        RECT  5.625 1.530 6.415 1.760 ;
        RECT  5.860 2.800 6.415 3.030 ;
        RECT  5.165 1.990 6.170 2.330 ;
        RECT  5.520 2.800 5.860 3.140 ;
        RECT  5.395 0.840 5.625 1.760 ;
        RECT  5.220 0.840 5.395 1.070 ;
        RECT  4.880 0.635 5.220 1.070 ;
        RECT  4.935 1.440 5.165 3.315 ;
        RECT  3.550 3.085 4.935 3.315 ;
        RECT  4.090 0.635 4.880 0.865 ;
        RECT  4.540 2.445 4.650 2.785 ;
        RECT  4.310 2.125 4.540 2.785 ;
        RECT  2.830 2.125 4.310 2.355 ;
        RECT  3.320 2.590 3.550 3.315 ;
        RECT  3.210 2.590 3.320 2.930 ;
        RECT  2.825 0.815 2.830 3.115 ;
        RECT  2.600 0.760 2.825 3.115 ;
        RECT  2.480 3.545 2.820 4.060 ;
        RECT  2.485 0.760 2.600 1.100 ;
        RECT  2.540 2.885 2.600 3.115 ;
        RECT  2.200 2.885 2.540 3.225 ;
        RECT  0.980 3.545 2.480 3.775 ;
        RECT  2.030 1.725 2.370 2.065 ;
        RECT  0.980 1.780 2.030 2.010 ;
        RECT  0.750 1.780 0.980 3.775 ;
        RECT  0.525 1.780 0.750 2.010 ;
        RECT  0.550 3.450 0.750 3.775 ;
        RECT  0.210 3.450 0.550 3.790 ;
        RECT  0.295 1.190 0.525 2.010 ;
        RECT  0.185 1.190 0.295 1.530 ;
    END
END DFFSX2

MACRO DFFSX1
    CLASS CORE ;
    FOREIGN DFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 3.900 9.790 4.410 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.460 0.870 11.690 3.870 ;
        RECT  10.945 0.870 11.460 1.100 ;
        RECT  11.100 3.640 11.460 3.870 ;
        RECT  10.760 3.640 11.100 4.370 ;
        RECT  10.605 0.670 10.945 1.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.325 2.630 12.360 3.210 ;
        RECT  12.095 1.250 12.325 3.210 ;
        RECT  11.960 1.250 12.095 1.590 ;
        RECT  12.020 2.630 12.095 3.210 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.080 1.845 1.580 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 2.965 1.105 3.195 ;
        RECT  0.725 2.575 0.955 3.195 ;
        RECT  0.555 2.575 0.725 2.805 ;
        RECT  0.215 2.465 0.555 2.805 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.685 -0.400 12.540 0.400 ;
        RECT  11.345 -0.400 11.685 0.575 ;
        RECT  10.220 -0.400 11.345 0.400 ;
        RECT  9.880 -0.400 10.220 0.960 ;
        RECT  8.560 -0.400 9.880 0.400 ;
        RECT  8.220 -0.400 8.560 0.575 ;
        RECT  6.165 -0.400 8.220 0.400 ;
        RECT  5.935 -0.400 6.165 1.010 ;
        RECT  4.040 -0.400 5.935 0.400 ;
        RECT  3.700 -0.400 4.040 1.110 ;
        RECT  1.545 -0.400 3.700 0.400 ;
        RECT  1.205 -0.400 1.545 0.575 ;
        RECT  0.000 -0.400 1.205 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 4.640 12.540 5.440 ;
        RECT  12.305 4.465 12.360 5.440 ;
        RECT  12.075 4.410 12.305 5.440 ;
        RECT  12.020 4.465 12.075 5.440 ;
        RECT  10.380 4.640 12.020 5.440 ;
        RECT  10.040 2.940 10.380 5.440 ;
        RECT  8.930 4.640 10.040 5.440 ;
        RECT  8.590 4.140 8.930 5.440 ;
        RECT  6.420 4.640 8.590 5.440 ;
        RECT  6.080 4.140 6.420 5.440 ;
        RECT  5.160 4.640 6.080 5.440 ;
        RECT  4.820 4.140 5.160 5.440 ;
        RECT  3.760 4.640 4.820 5.440 ;
        RECT  3.420 4.465 3.760 5.440 ;
        RECT  1.300 4.640 3.420 5.440 ;
        RECT  0.960 4.465 1.300 5.440 ;
        RECT  0.000 4.640 0.960 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.995 1.570 11.225 3.280 ;
        RECT  10.985 1.570 10.995 1.800 ;
        RECT  10.815 2.940 10.995 3.280 ;
        RECT  10.645 1.460 10.985 1.800 ;
        RECT  9.660 2.040 10.370 2.270 ;
        RECT  9.430 1.520 9.660 3.400 ;
        RECT  8.900 1.520 9.430 1.750 ;
        RECT  9.320 3.060 9.430 3.400 ;
        RECT  7.740 2.465 9.200 2.695 ;
        RECT  8.560 1.405 8.900 1.750 ;
        RECT  8.220 1.405 8.560 1.645 ;
        RECT  7.880 1.305 8.220 1.645 ;
        RECT  7.630 2.465 7.740 3.650 ;
        RECT  7.400 1.540 7.630 3.650 ;
        RECT  7.325 1.540 7.400 1.770 ;
        RECT  7.165 4.020 7.370 4.360 ;
        RECT  7.095 1.430 7.325 1.770 ;
        RECT  6.935 3.670 7.165 4.360 ;
        RECT  6.840 2.335 7.100 2.675 ;
        RECT  2.880 3.670 6.935 3.900 ;
        RECT  6.610 1.240 6.840 3.310 ;
        RECT  5.705 1.240 6.610 1.470 ;
        RECT  5.865 3.080 6.610 3.310 ;
        RECT  5.245 2.165 6.375 2.505 ;
        RECT  5.635 3.080 5.865 3.420 ;
        RECT  5.475 0.780 5.705 1.470 ;
        RECT  5.385 0.780 5.475 1.010 ;
        RECT  5.380 0.675 5.385 1.010 ;
        RECT  5.040 0.670 5.380 1.010 ;
        RECT  5.015 1.420 5.245 3.230 ;
        RECT  4.270 0.675 5.040 0.905 ;
        RECT  4.560 3.000 5.015 3.230 ;
        RECT  4.725 2.395 4.730 2.735 ;
        RECT  4.390 2.180 4.725 2.735 ;
        RECT  4.220 3.000 4.560 3.340 ;
        RECT  2.910 2.180 4.390 2.410 ;
        RECT  3.600 3.000 4.220 3.230 ;
        RECT  3.370 2.640 3.600 3.230 ;
        RECT  3.260 2.640 3.370 2.980 ;
        RECT  2.680 0.740 2.910 3.115 ;
        RECT  2.540 3.560 2.880 4.140 ;
        RECT  2.565 0.740 2.680 1.080 ;
        RECT  2.600 2.885 2.680 3.115 ;
        RECT  2.260 2.885 2.600 3.225 ;
        RECT  1.905 3.560 2.540 3.790 ;
        RECT  2.105 1.820 2.445 2.160 ;
        RECT  1.905 1.930 2.105 2.160 ;
        RECT  1.655 1.930 1.905 3.790 ;
        RECT  0.530 1.930 1.655 2.160 ;
        RECT  0.195 3.450 1.655 3.790 ;
        RECT  0.300 1.190 0.530 2.160 ;
        RECT  0.190 1.190 0.300 1.530 ;
    END
END DFFSX1

MACRO DFFRHQXL
    CLASS CORE ;
    FOREIGN DFFRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.610 2.910 12.400 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 3.715 13.660 4.055 ;
        RECT  13.415 1.305 13.645 4.055 ;
        RECT  12.755 1.305 13.415 1.535 ;
        RECT  13.320 3.715 13.415 4.055 ;
        RECT  12.650 1.260 12.755 1.535 ;
        RECT  12.310 1.195 12.650 1.535 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 1.680 1.840 2.110 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.170 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.870 -0.400 13.860 0.400 ;
        RECT  12.530 -0.400 12.870 0.575 ;
        RECT  11.365 -0.400 12.530 0.400 ;
        RECT  11.025 -0.400 11.365 0.575 ;
        RECT  9.765 -0.400 11.025 0.400 ;
        RECT  9.425 -0.400 9.765 0.575 ;
        RECT  6.790 -0.400 9.425 0.400 ;
        RECT  6.450 -0.400 6.790 1.160 ;
        RECT  4.100 -0.400 6.450 0.400 ;
        RECT  5.400 1.470 5.510 1.810 ;
        RECT  5.170 1.205 5.400 1.810 ;
        RECT  4.100 1.205 5.170 1.435 ;
        RECT  3.760 -0.400 4.100 1.435 ;
        RECT  1.480 -0.400 3.760 0.400 ;
        RECT  1.140 -0.400 1.480 0.575 ;
        RECT  0.000 -0.400 1.140 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.380 4.640 13.860 5.440 ;
        RECT  12.040 3.490 12.380 5.440 ;
        RECT  11.280 3.490 12.040 3.720 ;
        RECT  10.090 4.640 12.040 5.440 ;
        RECT  11.050 3.205 11.280 3.720 ;
        RECT  10.940 3.205 11.050 3.545 ;
        RECT  9.675 4.465 10.090 5.440 ;
        RECT  7.135 4.640 9.675 5.440 ;
        RECT  6.795 4.465 7.135 5.440 ;
        RECT  4.040 4.640 6.795 5.440 ;
        RECT  3.700 4.000 4.040 5.440 ;
        RECT  1.480 4.640 3.700 5.440 ;
        RECT  1.140 3.885 1.480 5.440 ;
        RECT  0.000 4.640 1.140 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.800 1.780 13.180 2.010 ;
        RECT  11.245 2.450 12.690 2.680 ;
        RECT  11.570 0.855 11.800 2.010 ;
        RECT  11.240 3.980 11.580 4.320 ;
        RECT  10.125 0.855 11.570 1.085 ;
        RECT  10.905 1.315 11.245 2.680 ;
        RECT  10.625 3.980 11.240 4.210 ;
        RECT  10.625 2.210 10.905 2.680 ;
        RECT  10.585 2.210 10.625 4.210 ;
        RECT  10.395 2.405 10.585 4.210 ;
        RECT  9.960 1.465 10.440 1.695 ;
        RECT  5.785 3.945 10.395 4.175 ;
        RECT  9.755 0.855 10.125 1.235 ;
        RECT  9.730 1.465 9.960 3.550 ;
        RECT  9.225 1.005 9.755 1.235 ;
        RECT  9.620 2.580 9.730 3.550 ;
        RECT  9.455 2.580 9.620 2.930 ;
        RECT  8.995 1.005 9.225 3.600 ;
        RECT  8.400 1.005 8.995 1.255 ;
        RECT  8.670 3.370 8.995 3.600 ;
        RECT  8.480 1.610 8.715 1.950 ;
        RECT  8.330 3.370 8.670 3.710 ;
        RECT  8.250 1.610 8.480 3.055 ;
        RECT  8.060 1.005 8.400 1.365 ;
        RECT  7.795 1.595 8.020 3.710 ;
        RECT  7.790 1.010 7.795 3.710 ;
        RECT  7.565 1.010 7.790 1.825 ;
        RECT  7.610 3.370 7.790 3.710 ;
        RECT  7.260 1.010 7.565 1.350 ;
        RECT  7.335 2.280 7.560 2.620 ;
        RECT  7.105 1.630 7.335 3.580 ;
        RECT  6.340 1.630 7.105 1.860 ;
        RECT  6.630 3.350 7.105 3.580 ;
        RECT  6.635 2.175 6.865 2.915 ;
        RECT  4.815 2.175 6.635 2.405 ;
        RECT  6.290 3.350 6.630 3.690 ;
        RECT  6.205 1.520 6.340 1.860 ;
        RECT  5.975 0.685 6.205 1.860 ;
        RECT  4.700 0.685 5.975 0.915 ;
        RECT  5.555 2.635 5.785 4.175 ;
        RECT  5.325 2.635 5.555 2.975 ;
        RECT  4.585 1.670 4.815 3.680 ;
        RECT  4.360 0.630 4.700 0.970 ;
        RECT  4.370 1.670 4.585 2.010 ;
        RECT  4.410 3.340 4.585 3.680 ;
        RECT  3.695 1.780 4.370 2.010 ;
        RECT  4.120 2.580 4.350 2.945 ;
        RECT  2.935 2.715 4.120 2.945 ;
        RECT  3.465 1.780 3.695 2.370 ;
        RECT  3.355 2.030 3.465 2.370 ;
        RECT  2.830 3.740 3.170 4.080 ;
        RECT  2.760 1.240 2.935 2.945 ;
        RECT  2.300 3.740 2.830 3.970 ;
        RECT  2.705 1.240 2.760 3.325 ;
        RECT  2.700 1.240 2.705 1.470 ;
        RECT  2.530 2.715 2.705 3.325 ;
        RECT  2.360 1.130 2.700 1.470 ;
        RECT  2.300 1.810 2.465 2.150 ;
        RECT  2.070 1.810 2.300 3.970 ;
        RECT  0.830 3.000 2.070 3.230 ;
        RECT  0.490 2.890 0.830 3.230 ;
        RECT  0.400 1.340 0.625 1.710 ;
        RECT  0.400 2.890 0.490 3.120 ;
        RECT  0.170 1.340 0.400 3.120 ;
    END
END DFFRHQXL

MACRO DFFRHQX4
    CLASS CORE ;
    FOREIGN DFFRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRHQXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.485 1.820 14.965 2.100 ;
        RECT  14.145 1.780 14.485 2.120 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.525 2.965 20.865 3.835 ;
        RECT  20.320 2.965 20.525 3.220 ;
        RECT  19.940 1.415 20.320 3.220 ;
        RECT  19.500 1.415 19.940 1.645 ;
        RECT  18.305 2.990 19.940 3.220 ;
        RECT  19.160 0.785 19.500 1.645 ;
        RECT  18.060 1.415 19.160 1.645 ;
        RECT  17.965 2.990 18.305 3.835 ;
        RECT  17.720 0.785 18.060 1.645 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.240 2.075 1.470 2.660 ;
        RECT  0.800 2.380 1.240 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.785 0.855 2.105 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.260 -0.400 21.120 0.400 ;
        RECT  19.920 -0.400 20.260 1.100 ;
        RECT  18.780 -0.400 19.920 0.400 ;
        RECT  18.440 -0.400 18.780 1.185 ;
        RECT  17.325 -0.400 18.440 0.400 ;
        RECT  16.985 -0.400 17.325 1.565 ;
        RECT  15.485 -0.400 16.985 0.400 ;
        RECT  15.145 -0.400 15.485 0.575 ;
        RECT  14.005 -0.400 15.145 0.400 ;
        RECT  13.665 -0.400 14.005 1.320 ;
        RECT  8.465 -0.400 13.665 0.400 ;
        RECT  8.125 -0.400 8.465 1.320 ;
        RECT  7.025 -0.400 8.125 0.400 ;
        RECT  6.685 -0.400 7.025 1.490 ;
        RECT  5.365 -0.400 6.685 0.400 ;
        RECT  5.365 1.260 5.405 1.600 ;
        RECT  5.065 -0.400 5.365 1.600 ;
        RECT  3.925 -0.400 5.065 0.400 ;
        RECT  3.585 -0.400 3.925 0.970 ;
        RECT  1.310 -0.400 3.585 0.400 ;
        RECT  0.970 -0.400 1.310 0.575 ;
        RECT  0.000 -0.400 0.970 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.585 4.640 21.120 5.440 ;
        RECT  19.245 3.450 19.585 5.440 ;
        RECT  16.970 4.640 19.245 5.440 ;
        RECT  16.740 3.110 16.970 5.440 ;
        RECT  15.325 4.640 16.740 5.440 ;
        RECT  14.985 4.465 15.325 5.440 ;
        RECT  13.625 4.640 14.985 5.440 ;
        RECT  13.395 4.080 13.625 5.440 ;
        RECT  8.685 4.640 13.395 5.440 ;
        RECT  8.345 4.465 8.685 5.440 ;
        RECT  7.160 4.640 8.345 5.440 ;
        RECT  6.930 4.040 7.160 5.440 ;
        RECT  5.735 4.640 6.930 5.440 ;
        RECT  5.395 4.465 5.735 5.440 ;
        RECT  3.845 4.640 5.395 5.440 ;
        RECT  3.505 4.465 3.845 5.440 ;
        RECT  1.200 4.640 3.505 5.440 ;
        RECT  1.200 3.485 1.255 3.825 ;
        RECT  0.970 3.485 1.200 5.440 ;
        RECT  0.915 3.485 0.970 3.825 ;
        RECT  0.000 4.640 0.970 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.880 2.045 19.220 2.385 ;
        RECT  16.785 2.125 18.880 2.355 ;
        RECT  16.755 2.125 16.785 2.550 ;
        RECT  16.525 0.805 16.755 2.550 ;
        RECT  14.725 0.805 16.525 1.035 ;
        RECT  16.510 2.125 16.525 2.550 ;
        RECT  16.280 2.125 16.510 4.140 ;
        RECT  16.065 1.265 16.295 1.605 ;
        RECT  14.490 3.910 16.280 4.140 ;
        RECT  15.565 1.375 16.065 1.605 ;
        RECT  15.820 2.200 16.050 3.570 ;
        RECT  14.660 3.340 15.820 3.570 ;
        RECT  15.335 1.375 15.565 3.110 ;
        RECT  13.745 2.360 15.335 2.590 ;
        RECT  14.385 0.805 14.725 1.330 ;
        RECT  14.430 3.160 14.660 3.570 ;
        RECT  14.150 3.910 14.490 4.250 ;
        RECT  13.135 3.160 14.430 3.390 ;
        RECT  13.920 3.620 14.150 4.140 ;
        RECT  13.160 3.620 13.920 3.850 ;
        RECT  13.515 2.245 13.745 2.590 ;
        RECT  13.265 2.245 13.515 2.475 ;
        RECT  12.925 2.135 13.265 2.475 ;
        RECT  12.930 3.620 13.160 4.365 ;
        RECT  12.905 2.780 13.135 3.390 ;
        RECT  9.145 4.135 12.930 4.365 ;
        RECT  12.510 2.780 12.905 3.010 ;
        RECT  12.615 3.280 12.670 3.620 ;
        RECT  12.510 1.100 12.645 1.440 ;
        RECT  12.330 3.280 12.615 3.845 ;
        RECT  12.280 0.675 12.510 3.010 ;
        RECT  9.725 3.615 12.330 3.845 ;
        RECT  11.205 0.675 12.280 0.905 ;
        RECT  12.055 2.635 12.280 3.010 ;
        RECT  10.820 2.635 12.055 2.865 ;
        RECT  11.815 1.140 11.925 1.480 ;
        RECT  11.585 1.140 11.815 1.840 ;
        RECT  10.485 1.610 11.585 1.840 ;
        RECT  10.185 3.095 11.580 3.325 ;
        RECT  10.865 0.675 11.205 1.380 ;
        RECT  9.385 0.675 10.865 0.905 ;
        RECT  10.535 2.520 10.820 2.865 ;
        RECT  10.480 2.520 10.535 2.860 ;
        RECT  10.145 1.140 10.485 1.840 ;
        RECT  10.120 2.905 10.185 3.325 ;
        RECT  10.120 1.310 10.145 1.840 ;
        RECT  9.955 1.310 10.120 3.325 ;
        RECT  9.890 1.310 9.955 3.190 ;
        RECT  9.185 1.310 9.890 1.540 ;
        RECT  9.715 2.850 9.890 3.190 ;
        RECT  9.495 3.425 9.725 3.845 ;
        RECT  8.650 2.905 9.715 3.135 ;
        RECT  9.430 1.770 9.660 2.435 ;
        RECT  8.080 3.425 9.495 3.655 ;
        RECT  8.080 2.205 9.430 2.435 ;
        RECT  8.845 1.310 9.185 1.785 ;
        RECT  8.915 4.005 9.145 4.365 ;
        RECT  7.620 4.005 8.915 4.235 ;
        RECT  7.745 1.555 8.845 1.785 ;
        RECT  8.310 2.770 8.650 3.135 ;
        RECT  7.850 2.205 8.080 3.655 ;
        RECT  7.150 2.205 7.850 2.435 ;
        RECT  7.515 1.150 7.745 1.785 ;
        RECT  7.390 3.295 7.620 4.235 ;
        RECT  7.405 1.150 7.515 1.490 ;
        RECT  6.535 3.295 7.390 3.525 ;
        RECT  7.095 2.205 7.150 3.060 ;
        RECT  6.865 1.775 7.095 3.060 ;
        RECT  6.300 1.775 6.865 2.005 ;
        RECT  6.810 2.720 6.865 3.060 ;
        RECT  6.400 3.880 6.630 4.225 ;
        RECT  6.305 2.235 6.535 3.525 ;
        RECT  3.040 3.995 6.400 4.225 ;
        RECT  5.335 2.235 6.305 2.465 ;
        RECT  6.190 1.260 6.300 2.005 ;
        RECT  5.960 0.675 6.190 2.005 ;
        RECT  5.735 2.930 6.075 3.300 ;
        RECT  5.595 0.675 5.960 0.905 ;
        RECT  4.765 2.930 5.735 3.160 ;
        RECT  4.995 2.110 5.335 2.465 ;
        RECT  4.535 1.140 4.765 3.160 ;
        RECT  4.345 1.140 4.535 1.480 ;
        RECT  4.380 2.930 4.535 3.160 ;
        RECT  4.040 2.930 4.380 3.270 ;
        RECT  3.945 2.040 4.285 2.640 ;
        RECT  3.615 2.930 4.040 3.160 ;
        RECT  2.735 2.040 3.945 2.270 ;
        RECT  3.275 2.570 3.615 3.160 ;
        RECT  2.810 2.670 3.040 4.225 ;
        RECT  2.645 2.670 2.810 3.065 ;
        RECT  1.950 3.995 2.810 4.225 ;
        RECT  2.505 0.900 2.735 2.270 ;
        RECT  2.415 3.420 2.550 3.760 ;
        RECT  2.305 0.900 2.505 1.240 ;
        RECT  2.415 2.040 2.505 2.270 ;
        RECT  2.185 2.040 2.415 3.760 ;
        RECT  1.950 1.470 2.275 1.810 ;
        RECT  1.720 1.275 1.950 4.225 ;
        RECT  0.535 1.275 1.720 1.505 ;
        RECT  0.535 2.890 1.720 3.245 ;
        RECT  0.195 0.695 0.535 1.505 ;
        RECT  0.195 2.890 0.535 4.170 ;
    END
END DFFRHQX4

MACRO DFFRHQX2
    CLASS CORE ;
    FOREIGN DFFRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRHQXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.415 2.655 13.950 3.205 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.160 1.210 16.390 3.105 ;
        RECT  15.030 1.210 16.160 1.440 ;
        RECT  15.700 2.875 16.160 3.105 ;
        RECT  15.360 2.875 15.700 4.030 ;
        RECT  14.690 0.635 15.030 1.445 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.645 1.720 1.840 2.085 ;
        RECT  1.280 1.720 1.645 2.140 ;
        RECT  1.250 1.720 1.280 2.085 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.020 2.380 1.105 2.635 ;
        RECT  0.600 2.230 1.020 2.680 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.790 -0.400 17.160 0.400 ;
        RECT  15.450 -0.400 15.790 0.575 ;
        RECT  14.045 -0.400 15.450 0.400 ;
        RECT  13.105 -0.400 14.045 0.575 ;
        RECT  11.760 -0.400 13.105 0.400 ;
        RECT  11.420 -0.400 11.760 0.575 ;
        RECT  7.845 -0.400 11.420 0.400 ;
        RECT  7.505 -0.400 7.845 1.290 ;
        RECT  3.950 -0.400 7.505 0.400 ;
        RECT  5.340 1.435 5.450 1.775 ;
        RECT  5.110 1.205 5.340 1.775 ;
        RECT  3.950 1.205 5.110 1.435 ;
        RECT  3.610 -0.400 3.950 1.435 ;
        RECT  1.325 -0.400 3.610 0.400 ;
        RECT  0.985 -0.400 1.325 0.575 ;
        RECT  0.000 -0.400 0.985 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.980 4.640 17.160 5.440 ;
        RECT  16.640 3.295 16.980 5.440 ;
        RECT  14.330 4.640 16.640 5.440 ;
        RECT  13.990 4.465 14.330 5.440 ;
        RECT  12.930 4.640 13.990 5.440 ;
        RECT  12.590 4.465 12.930 5.440 ;
        RECT  11.745 4.640 12.590 5.440 ;
        RECT  11.305 4.465 11.745 5.440 ;
        RECT  7.865 4.640 11.305 5.440 ;
        RECT  7.525 4.465 7.865 5.440 ;
        RECT  4.040 4.640 7.525 5.440 ;
        RECT  3.700 4.000 4.040 5.440 ;
        RECT  1.540 4.640 3.700 5.440 ;
        RECT  1.200 3.835 1.540 5.440 ;
        RECT  0.000 4.640 1.200 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.350 2.305 15.930 2.645 ;
        RECT  15.120 1.675 15.350 2.645 ;
        RECT  14.155 1.675 15.120 1.905 ;
        RECT  14.390 2.170 14.730 2.570 ;
        RECT  13.690 2.170 14.390 2.400 ;
        RECT  13.925 0.865 14.155 1.905 ;
        RECT  12.305 0.865 13.925 1.095 ;
        RECT  13.450 3.610 13.790 3.950 ;
        RECT  13.350 1.480 13.690 2.400 ;
        RECT  12.950 3.610 13.450 3.840 ;
        RECT  12.950 2.170 13.350 2.400 ;
        RECT  12.840 2.170 12.950 3.840 ;
        RECT  12.610 2.170 12.840 4.175 ;
        RECT  12.290 1.410 12.630 1.750 ;
        RECT  10.425 3.945 12.610 4.175 ;
        RECT  11.950 0.865 12.305 1.145 ;
        RECT  11.910 1.520 12.290 1.750 ;
        RECT  10.395 0.865 11.950 1.095 ;
        RECT  11.570 1.520 11.910 3.500 ;
        RECT  11.565 1.520 11.570 2.880 ;
        RECT  11.290 2.540 11.565 2.880 ;
        RECT  10.570 1.510 10.680 1.850 ;
        RECT  10.340 1.510 10.570 3.000 ;
        RECT  10.195 3.945 10.425 4.365 ;
        RECT  10.055 0.660 10.395 1.095 ;
        RECT  10.190 2.660 10.340 3.000 ;
        RECT  8.325 4.135 10.195 4.365 ;
        RECT  9.965 3.340 10.160 3.680 ;
        RECT  9.290 0.865 10.055 1.095 ;
        RECT  9.960 1.420 10.015 1.760 ;
        RECT  9.960 3.340 9.965 3.845 ;
        RECT  9.730 1.420 9.960 3.845 ;
        RECT  9.675 1.420 9.730 1.760 ;
        RECT  8.785 3.615 9.730 3.845 ;
        RECT  9.290 2.960 9.440 3.300 ;
        RECT  9.060 0.865 9.290 3.300 ;
        RECT  8.950 1.420 9.060 1.760 ;
        RECT  8.660 3.365 8.785 3.845 ;
        RECT  8.565 1.520 8.660 3.845 ;
        RECT  8.555 1.210 8.565 3.845 ;
        RECT  8.430 1.210 8.555 3.710 ;
        RECT  8.225 1.210 8.430 1.750 ;
        RECT  8.380 3.370 8.430 3.710 ;
        RECT  7.340 3.425 8.380 3.655 ;
        RECT  8.095 3.945 8.325 4.365 ;
        RECT  7.070 1.520 8.225 1.750 ;
        RECT  7.970 1.980 8.200 3.135 ;
        RECT  5.660 3.945 8.095 4.175 ;
        RECT  6.605 1.980 7.970 2.210 ;
        RECT  6.640 2.905 7.970 3.135 ;
        RECT  6.145 2.445 7.580 2.675 ;
        RECT  7.000 3.370 7.340 3.710 ;
        RECT  6.840 1.060 7.070 1.750 ;
        RECT  6.410 2.905 6.640 3.545 ;
        RECT  6.375 1.330 6.605 2.210 ;
        RECT  6.300 3.205 6.410 3.545 ;
        RECT  6.255 1.330 6.375 1.560 ;
        RECT  6.145 1.220 6.255 1.560 ;
        RECT  5.915 0.740 6.145 1.560 ;
        RECT  5.915 2.005 6.145 2.675 ;
        RECT  4.600 0.740 5.915 0.970 ;
        RECT  4.795 2.005 5.915 2.235 ;
        RECT  5.660 2.550 5.665 2.890 ;
        RECT  5.430 2.550 5.660 4.175 ;
        RECT  5.325 2.550 5.430 2.890 ;
        RECT  4.650 1.780 4.795 3.680 ;
        RECT  4.565 1.670 4.650 3.680 ;
        RECT  4.260 0.630 4.600 0.970 ;
        RECT  4.310 1.670 4.565 2.010 ;
        RECT  4.415 3.340 4.565 3.680 ;
        RECT  3.995 2.550 4.335 2.945 ;
        RECT  3.665 1.780 4.310 2.010 ;
        RECT  2.895 2.715 3.995 2.945 ;
        RECT  3.435 1.780 3.665 2.480 ;
        RECT  3.325 2.140 3.435 2.480 ;
        RECT  3.050 3.790 3.105 4.130 ;
        RECT  2.765 3.785 3.050 4.130 ;
        RECT  2.665 1.395 2.895 3.325 ;
        RECT  2.305 3.785 2.765 4.015 ;
        RECT  2.585 1.395 2.665 1.625 ;
        RECT  2.535 2.930 2.665 3.325 ;
        RECT  2.245 0.815 2.585 1.625 ;
        RECT  2.075 1.855 2.305 4.015 ;
        RECT  0.780 2.910 2.075 3.140 ;
        RECT  0.440 2.910 0.780 3.720 ;
        RECT  0.360 1.195 0.665 1.535 ;
        RECT  0.360 2.910 0.440 3.140 ;
        RECT  0.130 1.195 0.360 3.140 ;
    END
END DFFRHQX2

MACRO DFFRHQX1
    CLASS CORE ;
    FOREIGN DFFRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRHQXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.610 2.910 12.400 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.630 1.245 13.645 3.195 ;
        RECT  13.415 1.245 13.630 4.290 ;
        RECT  12.570 1.245 13.415 1.475 ;
        RECT  13.340 2.965 13.415 4.290 ;
        RECT  13.290 3.480 13.340 4.290 ;
        RECT  12.340 0.730 12.570 1.475 ;
        RECT  12.230 0.730 12.340 1.070 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.615 1.285 1.765 1.515 ;
        RECT  1.615 1.810 1.620 2.150 ;
        RECT  1.385 1.285 1.615 2.150 ;
        RECT  1.280 1.810 1.385 2.150 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 2.405 1.105 2.660 ;
        RECT  0.580 2.170 0.900 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.290 -0.400 13.860 0.400 ;
        RECT  12.950 -0.400 13.290 0.950 ;
        RECT  11.805 -0.400 12.950 0.400 ;
        RECT  10.865 -0.400 11.805 0.575 ;
        RECT  9.725 -0.400 10.865 0.400 ;
        RECT  9.385 -0.400 9.725 0.575 ;
        RECT  6.795 -0.400 9.385 0.400 ;
        RECT  6.455 -0.400 6.795 1.130 ;
        RECT  4.020 -0.400 6.455 0.400 ;
        RECT  5.360 1.480 5.470 1.820 ;
        RECT  5.130 1.205 5.360 1.820 ;
        RECT  4.020 1.205 5.130 1.435 ;
        RECT  3.680 -0.400 4.020 1.435 ;
        RECT  1.295 -0.400 3.680 0.400 ;
        RECT  0.955 -0.400 1.295 1.045 ;
        RECT  0.000 -0.400 0.955 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.350 4.640 13.860 5.440 ;
        RECT  12.010 3.520 12.350 5.440 ;
        RECT  11.280 3.535 12.010 3.765 ;
        RECT  10.090 4.640 12.010 5.440 ;
        RECT  11.050 2.930 11.280 3.765 ;
        RECT  10.940 2.930 11.050 3.270 ;
        RECT  9.675 4.465 10.090 5.440 ;
        RECT  7.215 4.640 9.675 5.440 ;
        RECT  6.800 4.465 7.215 5.440 ;
        RECT  4.040 4.640 6.800 5.440 ;
        RECT  3.700 3.980 4.040 5.440 ;
        RECT  1.580 4.640 3.700 5.440 ;
        RECT  1.240 3.800 1.580 5.440 ;
        RECT  0.000 4.640 1.240 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.810 1.710 13.150 2.050 ;
        RECT  11.760 1.710 12.810 1.940 ;
        RECT  11.240 2.450 12.690 2.680 ;
        RECT  11.530 0.865 11.760 1.940 ;
        RECT  11.285 4.000 11.625 4.340 ;
        RECT  10.085 0.865 11.530 1.095 ;
        RECT  10.705 4.000 11.285 4.230 ;
        RECT  10.925 1.375 11.240 2.680 ;
        RECT  10.865 1.375 10.925 1.715 ;
        RECT  10.705 2.210 10.925 2.680 ;
        RECT  10.585 2.210 10.705 4.230 ;
        RECT  10.475 2.405 10.585 4.230 ;
        RECT  10.470 3.945 10.475 4.230 ;
        RECT  5.785 3.945 10.470 4.175 ;
        RECT  10.060 1.410 10.400 1.750 ;
        RECT  9.715 0.865 10.085 1.145 ;
        RECT  10.040 1.520 10.060 1.750 ;
        RECT  9.810 1.520 10.040 3.500 ;
        RECT  9.620 2.580 9.810 3.500 ;
        RECT  9.225 0.865 9.715 1.095 ;
        RECT  9.455 2.580 9.620 2.930 ;
        RECT  8.995 0.865 9.225 3.600 ;
        RECT  8.305 0.865 8.995 1.105 ;
        RECT  8.670 3.370 8.995 3.600 ;
        RECT  8.480 1.605 8.675 1.945 ;
        RECT  8.330 3.370 8.670 3.710 ;
        RECT  8.335 1.605 8.480 3.055 ;
        RECT  8.250 1.610 8.335 3.055 ;
        RECT  8.075 0.865 8.305 1.275 ;
        RECT  7.950 1.595 8.020 3.705 ;
        RECT  7.815 1.595 7.950 3.710 ;
        RECT  7.790 1.120 7.815 3.710 ;
        RECT  7.585 1.120 7.790 1.825 ;
        RECT  7.610 3.370 7.790 3.710 ;
        RECT  7.560 1.120 7.585 1.350 ;
        RECT  7.220 1.010 7.560 1.350 ;
        RECT  7.335 2.300 7.560 2.705 ;
        RECT  7.105 1.640 7.335 3.580 ;
        RECT  6.300 1.640 7.105 1.870 ;
        RECT  6.630 3.350 7.105 3.580 ;
        RECT  6.635 2.175 6.865 2.915 ;
        RECT  4.865 2.175 6.635 2.405 ;
        RECT  6.290 3.350 6.630 3.690 ;
        RECT  6.165 1.530 6.300 1.870 ;
        RECT  5.935 0.740 6.165 1.870 ;
        RECT  4.660 0.740 5.935 0.970 ;
        RECT  5.555 2.635 5.785 4.175 ;
        RECT  5.320 2.635 5.555 2.975 ;
        RECT  4.670 1.780 4.865 3.680 ;
        RECT  4.635 1.670 4.670 3.680 ;
        RECT  4.320 0.630 4.660 0.970 ;
        RECT  4.330 1.670 4.635 2.010 ;
        RECT  4.410 3.340 4.635 3.680 ;
        RECT  4.065 2.580 4.405 2.945 ;
        RECT  3.630 1.780 4.330 2.010 ;
        RECT  2.895 2.715 4.065 2.945 ;
        RECT  3.400 1.780 3.630 2.370 ;
        RECT  3.290 2.030 3.400 2.370 ;
        RECT  2.830 3.740 3.170 4.080 ;
        RECT  2.850 1.045 2.895 2.945 ;
        RECT  2.665 1.045 2.850 3.325 ;
        RECT  2.280 3.740 2.830 3.970 ;
        RECT  2.660 1.045 2.665 1.275 ;
        RECT  2.615 2.715 2.665 3.325 ;
        RECT  2.320 0.935 2.660 1.275 ;
        RECT  2.510 2.985 2.615 3.325 ;
        RECT  2.280 1.830 2.335 2.170 ;
        RECT  2.050 1.830 2.280 3.970 ;
        RECT  1.995 1.830 2.050 2.170 ;
        RECT  0.780 2.890 2.050 3.120 ;
        RECT  0.440 2.890 0.780 3.230 ;
        RECT  0.350 1.280 0.520 1.620 ;
        RECT  0.350 2.890 0.440 3.120 ;
        RECT  0.120 1.280 0.350 3.120 ;
    END
END DFFRHQX1

MACRO DFFRXL
    CLASS CORE ;
    FOREIGN DFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 2.860 4.480 3.280 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.010 0.865 14.240 3.755 ;
        RECT  13.410 0.865 14.010 1.095 ;
        RECT  13.695 3.525 14.010 3.755 ;
        RECT  13.645 3.525 13.695 4.035 ;
        RECT  13.315 3.500 13.645 4.035 ;
        RECT  13.070 0.635 13.410 1.095 ;
        RECT  13.250 3.805 13.315 4.035 ;
        RECT  12.910 3.805 13.250 4.230 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.835 1.820 15.040 2.100 ;
        RECT  14.835 3.620 14.920 3.960 ;
        RECT  14.820 1.820 14.835 3.960 ;
        RECT  14.605 1.265 14.820 3.960 ;
        RECT  14.475 1.265 14.605 2.075 ;
        RECT  14.580 3.620 14.605 3.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.740 1.960 2.080 ;
        RECT  1.620 1.740 1.765 2.105 ;
        RECT  1.320 1.795 1.620 2.105 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.550 1.265 3.220 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 -0.400 15.180 0.400 ;
        RECT  13.800 -0.400 14.140 0.575 ;
        RECT  12.530 -0.400 13.800 0.400 ;
        RECT  12.190 -0.400 12.530 0.950 ;
        RECT  10.770 -0.400 12.190 0.400 ;
        RECT  10.430 -0.400 10.770 1.300 ;
        RECT  6.170 -0.400 10.430 0.400 ;
        RECT  7.870 1.420 7.880 1.760 ;
        RECT  7.540 1.205 7.870 1.760 ;
        RECT  6.580 1.205 7.540 1.435 ;
        RECT  6.240 1.205 6.580 1.560 ;
        RECT  6.170 1.205 6.240 1.505 ;
        RECT  5.940 -0.400 6.170 1.505 ;
        RECT  4.655 -0.400 5.940 0.400 ;
        RECT  4.315 -0.400 4.655 0.960 ;
        RECT  1.555 -0.400 4.315 0.400 ;
        RECT  1.215 -0.400 1.555 0.575 ;
        RECT  0.000 -0.400 1.215 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.150 4.640 15.180 5.440 ;
        RECT  13.810 4.465 14.150 5.440 ;
        RECT  12.530 4.640 13.810 5.440 ;
        RECT  12.190 4.085 12.530 5.440 ;
        RECT  10.465 4.640 12.190 5.440 ;
        RECT  10.125 4.080 10.465 5.440 ;
        RECT  8.370 4.640 10.125 5.440 ;
        RECT  7.430 4.080 8.370 5.440 ;
        RECT  4.070 4.640 7.430 5.440 ;
        RECT  3.730 4.465 4.070 5.440 ;
        RECT  1.480 4.640 3.730 5.440 ;
        RECT  1.140 4.465 1.480 5.440 ;
        RECT  0.000 4.640 1.140 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.495 1.545 13.725 3.105 ;
        RECT  13.355 1.545 13.495 1.775 ;
        RECT  13.085 2.875 13.495 3.105 ;
        RECT  13.125 1.420 13.355 1.775 ;
        RECT  12.440 2.110 13.100 2.450 ;
        RECT  12.855 2.875 13.085 3.350 ;
        RECT  12.210 1.865 12.440 3.760 ;
        RECT  11.650 1.865 12.210 2.095 ;
        RECT  11.170 3.530 12.210 3.760 ;
        RECT  11.285 0.915 11.650 2.095 ;
        RECT  10.240 3.060 11.535 3.290 ;
        RECT  10.930 1.865 11.285 2.095 ;
        RECT  10.830 3.530 11.170 3.960 ;
        RECT  10.830 1.865 10.930 2.570 ;
        RECT  10.700 1.865 10.830 2.580 ;
        RECT  10.490 2.240 10.700 2.580 ;
        RECT  10.010 1.550 10.240 3.290 ;
        RECT  9.315 1.550 10.010 1.780 ;
        RECT  9.765 3.060 10.010 3.290 ;
        RECT  9.465 3.060 9.765 4.340 ;
        RECT  9.240 2.390 9.470 2.790 ;
        RECT  9.425 4.000 9.465 4.340 ;
        RECT  9.085 1.290 9.315 1.780 ;
        RECT  8.875 2.560 9.240 2.790 ;
        RECT  8.645 2.560 8.875 3.850 ;
        RECT  8.415 2.090 8.855 2.320 ;
        RECT  7.185 3.620 8.645 3.850 ;
        RECT  8.185 0.675 8.415 3.385 ;
        RECT  6.745 0.675 8.185 0.905 ;
        RECT  7.430 3.155 8.185 3.385 ;
        RECT  7.685 2.305 7.915 2.670 ;
        RECT  6.725 2.305 7.685 2.560 ;
        RECT  6.955 2.810 7.185 4.365 ;
        RECT  4.530 4.135 6.955 4.365 ;
        RECT  6.405 0.635 6.745 0.975 ;
        RECT  6.495 1.825 6.725 3.690 ;
        RECT  5.705 1.825 6.495 2.055 ;
        RECT  5.750 3.460 6.495 3.690 ;
        RECT  5.925 2.440 6.265 2.780 ;
        RECT  5.015 2.495 5.925 2.725 ;
        RECT  5.410 3.460 5.750 3.800 ;
        RECT  5.475 1.100 5.705 2.055 ;
        RECT  3.875 1.655 5.475 1.885 ;
        RECT  5.120 0.770 5.230 1.110 ;
        RECT  4.890 0.770 5.120 1.420 ;
        RECT  4.990 2.115 5.015 2.725 ;
        RECT  4.760 2.115 4.990 3.870 ;
        RECT  3.305 1.190 4.890 1.420 ;
        RECT  4.675 2.115 4.760 2.455 ;
        RECT  4.300 4.005 4.530 4.365 ;
        RECT  3.345 4.005 4.300 4.235 ;
        RECT  3.535 1.655 3.875 2.080 ;
        RECT  3.115 4.005 3.345 4.320 ;
        RECT  3.075 1.190 3.305 3.605 ;
        RECT  2.325 4.090 3.115 4.320 ;
        RECT  2.915 1.190 3.075 1.420 ;
        RECT  2.785 3.375 3.075 3.605 ;
        RECT  2.575 0.965 2.915 1.420 ;
        RECT  2.555 3.375 2.785 3.800 ;
        RECT  2.350 1.890 2.580 3.060 ;
        RECT  2.325 2.830 2.350 3.060 ;
        RECT  2.095 2.830 2.325 4.320 ;
        RECT  2.075 3.995 2.095 4.320 ;
        RECT  0.765 3.995 2.075 4.225 ;
        RECT  0.600 1.110 0.940 1.450 ;
        RECT  0.545 3.515 0.765 4.225 ;
        RECT  0.545 1.220 0.600 1.450 ;
        RECT  0.315 1.220 0.545 4.225 ;
    END
END DFFRXL

MACRO DFFRX4
    CLASS CORE ;
    FOREIGN DFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 2.745 4.480 3.495 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.300 1.195 17.680 3.220 ;
        RECT  17.280 1.195 17.300 1.535 ;
        RECT  17.280 2.780 17.300 3.120 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.900 1.260 19.000 3.120 ;
        RECT  18.620 1.195 18.900 3.120 ;
        RECT  18.615 1.195 18.620 2.075 ;
        RECT  18.560 2.780 18.620 3.120 ;
        RECT  18.560 1.195 18.615 1.535 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 2.710 1.845 3.295 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 1.850 1.180 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.540 -0.400 19.800 0.400 ;
        RECT  19.200 -0.400 19.540 0.950 ;
        RECT  18.260 -0.400 19.200 0.400 ;
        RECT  17.920 -0.400 18.260 0.950 ;
        RECT  16.980 -0.400 17.920 0.400 ;
        RECT  16.640 -0.400 16.980 0.950 ;
        RECT  15.610 -0.400 16.640 0.400 ;
        RECT  15.270 -0.400 15.610 0.950 ;
        RECT  14.170 -0.400 15.270 0.400 ;
        RECT  13.830 -0.400 14.170 0.950 ;
        RECT  12.710 -0.400 13.830 0.400 ;
        RECT  12.370 -0.400 12.710 0.950 ;
        RECT  10.940 -0.400 12.370 0.400 ;
        RECT  10.600 -0.400 10.940 1.080 ;
        RECT  8.345 -0.400 10.600 0.400 ;
        RECT  8.115 -0.400 8.345 1.475 ;
        RECT  6.490 -0.400 8.115 0.400 ;
        RECT  7.930 1.245 8.115 1.475 ;
        RECT  6.150 -0.400 6.490 0.960 ;
        RECT  4.865 -0.400 6.150 0.400 ;
        RECT  4.525 -0.400 4.865 1.335 ;
        RECT  1.295 -0.400 4.525 0.400 ;
        RECT  0.955 -0.400 1.295 0.575 ;
        RECT  0.000 -0.400 0.955 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.540 4.640 19.800 5.440 ;
        RECT  19.200 4.040 19.540 5.440 ;
        RECT  18.260 4.640 19.200 5.440 ;
        RECT  17.920 4.040 18.260 5.440 ;
        RECT  16.980 4.640 17.920 5.440 ;
        RECT  16.640 4.040 16.980 5.440 ;
        RECT  15.410 4.640 16.640 5.440 ;
        RECT  15.070 2.845 15.410 5.440 ;
        RECT  12.810 4.640 15.070 5.440 ;
        RECT  12.470 4.080 12.810 5.440 ;
        RECT  10.330 4.640 12.470 5.440 ;
        RECT  9.990 3.675 10.330 5.440 ;
        RECT  7.480 4.640 9.990 5.440 ;
        RECT  7.140 3.920 7.480 5.440 ;
        RECT  3.820 4.640 7.140 5.440 ;
        RECT  3.480 4.465 3.820 5.440 ;
        RECT  1.545 4.640 3.480 5.440 ;
        RECT  1.150 4.385 1.545 5.440 ;
        RECT  0.000 4.640 1.150 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.305 2.030 19.535 3.750 ;
        RECT  16.975 3.520 19.305 3.750 ;
        RECT  16.745 1.395 16.975 3.750 ;
        RECT  16.290 1.395 16.745 1.730 ;
        RECT  16.130 3.265 16.745 3.495 ;
        RECT  15.510 2.100 16.450 2.440 ;
        RECT  15.950 1.390 16.290 1.730 ;
        RECT  15.790 2.975 16.130 3.785 ;
        RECT  15.940 1.395 15.950 1.675 ;
        RECT  14.890 2.155 15.510 2.385 ;
        RECT  14.660 0.720 14.890 2.690 ;
        RECT  14.550 0.720 14.660 1.475 ;
        RECT  14.130 2.460 14.660 2.690 ;
        RECT  13.450 1.245 14.550 1.475 ;
        RECT  14.055 1.725 14.410 2.065 ;
        RECT  13.900 2.460 14.130 3.835 ;
        RECT  13.470 1.725 14.055 2.105 ;
        RECT  13.790 2.985 13.900 3.835 ;
        RECT  12.200 3.605 13.790 3.835 ;
        RECT  12.465 1.875 13.470 2.105 ;
        RECT  13.220 0.700 13.450 1.475 ;
        RECT  13.110 0.700 13.220 1.040 ;
        RECT  12.235 1.495 12.465 3.365 ;
        RECT  9.895 1.495 12.235 1.735 ;
        RECT  11.605 3.135 12.235 3.365 ;
        RECT  11.970 3.605 12.200 4.250 ;
        RECT  11.465 2.425 11.805 2.820 ;
        RECT  11.605 3.750 11.660 4.090 ;
        RECT  11.375 3.135 11.605 4.090 ;
        RECT  9.435 2.425 11.465 2.655 ;
        RECT  9.695 3.135 11.375 3.365 ;
        RECT  11.320 3.750 11.375 4.090 ;
        RECT  9.665 1.105 9.895 1.735 ;
        RECT  9.465 3.135 9.695 3.855 ;
        RECT  9.250 1.105 9.665 1.335 ;
        RECT  9.050 3.625 9.465 3.855 ;
        RECT  9.205 1.750 9.435 2.655 ;
        RECT  8.920 2.425 9.205 2.655 ;
        RECT  8.710 3.625 9.050 3.990 ;
        RECT  8.690 1.745 8.920 3.145 ;
        RECT  7.465 1.745 8.690 1.975 ;
        RECT  8.245 2.915 8.690 3.145 ;
        RECT  6.875 2.235 8.460 2.465 ;
        RECT  8.240 2.915 8.245 3.945 ;
        RECT  8.015 2.915 8.240 4.000 ;
        RECT  7.900 3.660 8.015 4.000 ;
        RECT  7.505 2.840 7.670 3.180 ;
        RECT  7.275 2.840 7.505 3.660 ;
        RECT  7.235 0.675 7.465 1.975 ;
        RECT  6.745 3.430 7.275 3.660 ;
        RECT  6.740 0.675 7.235 0.905 ;
        RECT  6.645 1.565 6.875 3.145 ;
        RECT  6.515 3.430 6.745 4.365 ;
        RECT  5.930 1.565 6.645 1.795 ;
        RECT  6.200 2.915 6.645 3.145 ;
        RECT  4.365 4.135 6.515 4.365 ;
        RECT  5.860 2.915 6.200 3.870 ;
        RECT  5.830 2.100 6.170 2.440 ;
        RECT  5.590 1.430 5.930 1.795 ;
        RECT  5.015 2.155 5.830 2.385 ;
        RECT  3.550 1.565 5.590 1.795 ;
        RECT  5.015 3.560 5.070 3.900 ;
        RECT  4.785 2.025 5.015 3.900 ;
        RECT  4.270 2.025 4.785 2.255 ;
        RECT  4.730 3.560 4.785 3.900 ;
        RECT  4.135 3.945 4.365 4.365 ;
        RECT  2.575 0.825 4.275 1.055 ;
        RECT  3.165 3.945 4.135 4.175 ;
        RECT  3.550 2.320 3.660 2.660 ;
        RECT  3.320 1.565 3.550 2.660 ;
        RECT  2.955 3.035 3.165 4.400 ;
        RECT  2.935 1.775 2.955 4.400 ;
        RECT  2.725 1.775 2.935 3.265 ;
        RECT  2.020 4.170 2.935 4.400 ;
        RECT  2.090 1.775 2.725 2.005 ;
        RECT  2.490 3.500 2.620 3.840 ;
        RECT  2.345 0.825 2.575 1.470 ;
        RECT  2.260 2.240 2.490 3.840 ;
        RECT  2.235 1.130 2.345 1.470 ;
        RECT  1.850 2.240 2.260 2.470 ;
        RECT  1.850 1.185 2.235 1.415 ;
        RECT  1.790 3.710 2.020 4.400 ;
        RECT  1.620 1.185 1.850 2.470 ;
        RECT  0.605 3.710 1.790 3.940 ;
        RECT  0.495 1.220 0.635 1.560 ;
        RECT  0.495 3.010 0.605 3.940 ;
        RECT  0.295 1.220 0.495 3.940 ;
        RECT  0.265 1.275 0.295 3.940 ;
    END
END DFFRX4

MACRO DFFRX2
    CLASS CORE ;
    FOREIGN DFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.605 2.875 4.660 3.390 ;
        RECT  4.320 2.755 4.605 3.390 ;
        RECT  4.175 2.755 4.320 3.335 ;
        RECT  4.130 2.875 4.175 3.240 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.570 1.515 15.710 2.130 ;
        RECT  15.565 2.930 15.620 3.270 ;
        RECT  15.565 1.260 15.570 2.130 ;
        RECT  15.335 1.260 15.565 3.270 ;
        RECT  15.150 1.260 15.335 2.130 ;
        RECT  15.280 2.930 15.335 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.000 1.260 17.005 3.230 ;
        RECT  16.705 1.260 17.000 3.275 ;
        RECT  16.640 1.260 16.705 1.600 ;
        RECT  16.570 2.930 16.705 3.275 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.935 1.840 3.775 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.260 1.180 2.075 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.280 -0.400 17.160 0.400 ;
        RECT  15.940 -0.400 16.280 0.950 ;
        RECT  14.120 -0.400 15.940 0.400 ;
        RECT  13.780 -0.400 14.120 1.360 ;
        RECT  12.630 -0.400 13.780 0.400 ;
        RECT  12.290 -0.400 12.630 0.575 ;
        RECT  10.770 -0.400 12.290 0.400 ;
        RECT  10.430 -0.400 10.770 1.250 ;
        RECT  8.040 -0.400 10.430 0.400 ;
        RECT  7.700 -0.400 8.040 1.370 ;
        RECT  6.340 -0.400 7.700 0.400 ;
        RECT  6.000 -0.400 6.340 0.960 ;
        RECT  5.120 -0.400 6.000 0.440 ;
        RECT  4.695 -0.400 5.120 1.335 ;
        RECT  1.300 -0.400 4.695 0.400 ;
        RECT  0.960 -0.400 1.300 0.575 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.260 4.640 17.160 5.440 ;
        RECT  15.920 4.080 16.260 5.440 ;
        RECT  14.200 4.640 15.920 5.440 ;
        RECT  13.860 3.680 14.200 5.440 ;
        RECT  11.420 4.640 13.860 5.440 ;
        RECT  11.080 4.080 11.420 5.440 ;
        RECT  8.705 4.640 11.080 5.440 ;
        RECT  7.260 4.135 8.705 5.440 ;
        RECT  4.360 4.640 7.260 5.440 ;
        RECT  4.020 4.465 4.360 5.440 ;
        RECT  1.460 4.640 4.020 5.440 ;
        RECT  1.120 4.465 1.460 5.440 ;
        RECT  0.000 4.640 1.120 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.245 1.910 16.475 2.655 ;
        RECT  16.200 2.425 16.245 2.655 ;
        RECT  15.970 2.425 16.200 3.805 ;
        RECT  14.920 3.575 15.970 3.805 ;
        RECT  14.810 3.575 14.920 4.020 ;
        RECT  14.810 1.020 14.840 1.360 ;
        RECT  14.580 1.020 14.810 4.020 ;
        RECT  14.500 1.020 14.580 1.360 ;
        RECT  14.295 1.630 14.350 2.045 ;
        RECT  14.065 1.630 14.295 3.165 ;
        RECT  14.010 1.630 14.065 2.045 ;
        RECT  13.520 2.935 14.065 3.165 ;
        RECT  13.400 1.815 14.010 2.045 ;
        RECT  13.290 2.935 13.520 3.510 ;
        RECT  13.170 0.910 13.400 2.045 ;
        RECT  12.740 3.280 13.290 3.510 ;
        RECT  13.060 0.910 13.170 1.250 ;
        RECT  12.490 1.815 13.170 2.045 ;
        RECT  12.630 3.280 12.740 3.620 ;
        RECT  12.400 3.280 12.630 4.270 ;
        RECT  12.050 2.460 12.550 2.800 ;
        RECT  12.205 1.630 12.490 2.045 ;
        RECT  12.120 3.930 12.400 4.270 ;
        RECT  12.150 1.630 12.205 1.970 ;
        RECT  11.920 2.460 12.050 3.335 ;
        RECT  11.690 1.685 11.920 3.335 ;
        RECT  11.590 1.685 11.690 1.915 ;
        RECT  11.680 2.680 11.690 3.335 ;
        RECT  10.665 3.105 11.680 3.335 ;
        RECT  11.360 1.225 11.590 1.915 ;
        RECT  11.405 2.205 11.460 2.435 ;
        RECT  11.175 2.205 11.405 2.440 ;
        RECT  11.130 1.225 11.360 1.755 ;
        RECT  10.785 2.210 11.175 2.440 ;
        RECT  9.460 1.525 11.130 1.755 ;
        RECT  10.555 1.985 10.785 2.440 ;
        RECT  10.435 3.105 10.665 3.480 ;
        RECT  9.000 1.985 10.555 2.215 ;
        RECT  10.100 3.250 10.435 3.480 ;
        RECT  9.760 3.250 10.100 3.590 ;
        RECT  9.520 2.600 9.860 2.940 ;
        RECT  9.505 2.710 9.520 2.940 ;
        RECT  9.275 2.710 9.505 3.900 ;
        RECT  9.230 1.090 9.460 1.755 ;
        RECT  7.375 3.670 9.275 3.900 ;
        RECT  9.060 1.090 9.230 1.430 ;
        RECT  8.770 1.705 9.000 3.440 ;
        RECT  7.240 1.705 8.770 1.935 ;
        RECT  7.830 3.210 8.770 3.440 ;
        RECT  8.200 2.170 8.540 2.885 ;
        RECT  6.575 2.170 8.200 2.400 ;
        RECT  7.530 2.630 7.870 2.970 ;
        RECT  7.375 2.685 7.530 2.970 ;
        RECT  7.145 2.685 7.375 3.900 ;
        RECT  7.235 1.205 7.240 1.935 ;
        RECT  7.125 1.150 7.235 1.935 ;
        RECT  6.935 3.670 7.145 3.900 ;
        RECT  6.950 0.665 7.125 1.935 ;
        RECT  6.895 0.665 6.950 1.490 ;
        RECT  6.705 3.670 6.935 4.355 ;
        RECT  6.630 0.665 6.895 0.895 ;
        RECT  4.825 4.125 6.705 4.355 ;
        RECT  6.345 1.575 6.575 3.185 ;
        RECT  5.840 1.575 6.345 1.805 ;
        RECT  6.155 2.955 6.345 3.185 ;
        RECT  6.155 3.470 6.210 3.810 ;
        RECT  5.925 2.955 6.155 3.810 ;
        RECT  5.775 2.140 6.115 2.480 ;
        RECT  5.870 3.470 5.925 3.810 ;
        RECT  5.610 1.455 5.840 1.805 ;
        RECT  5.345 2.195 5.775 2.425 ;
        RECT  5.500 1.455 5.610 1.795 ;
        RECT  3.680 1.565 5.500 1.795 ;
        RECT  5.345 3.550 5.400 3.890 ;
        RECT  5.115 2.195 5.345 3.890 ;
        RECT  5.110 2.195 5.115 2.425 ;
        RECT  5.060 3.550 5.115 3.890 ;
        RECT  4.560 2.030 5.110 2.425 ;
        RECT  4.595 3.945 4.825 4.355 ;
        RECT  3.705 3.945 4.595 4.175 ;
        RECT  4.080 0.675 4.420 1.110 ;
        RECT  3.025 0.675 4.080 0.905 ;
        RECT  3.475 3.945 3.705 4.255 ;
        RECT  3.350 1.565 3.680 2.085 ;
        RECT  2.560 4.025 3.475 4.255 ;
        RECT  3.340 1.745 3.350 2.085 ;
        RECT  3.045 3.300 3.100 3.640 ;
        RECT  3.025 3.280 3.045 3.640 ;
        RECT  2.795 0.675 3.025 3.640 ;
        RECT  2.430 0.675 2.795 1.270 ;
        RECT  2.760 3.300 2.795 3.640 ;
        RECT  2.460 3.970 2.560 4.310 ;
        RECT  2.415 1.590 2.460 4.310 ;
        RECT  2.375 0.905 2.430 1.270 ;
        RECT  2.230 1.535 2.415 4.310 ;
        RECT  2.320 0.930 2.375 1.270 ;
        RECT  2.075 1.535 2.230 1.875 ;
        RECT  2.220 3.970 2.230 4.310 ;
        RECT  0.500 4.005 2.220 4.235 ;
        RECT  0.500 1.105 0.555 1.445 ;
        RECT  0.500 3.055 0.555 3.395 ;
        RECT  0.270 1.105 0.500 4.235 ;
        RECT  0.215 1.105 0.270 1.445 ;
        RECT  0.215 3.055 0.270 3.395 ;
    END
END DFFRX2

MACRO DFFRX1
    CLASS CORE ;
    FOREIGN DFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.525 3.340 4.825 3.570 ;
        RECT  4.130 2.950 4.525 3.570 ;
        RECT  4.100 2.965 4.130 3.570 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.180 2.035 14.410 3.295 ;
        RECT  13.575 2.035 14.180 2.265 ;
        RECT  13.890 3.065 14.180 3.295 ;
        RECT  13.660 3.065 13.890 3.795 ;
        RECT  13.520 3.500 13.660 3.795 ;
        RECT  13.345 1.380 13.575 2.265 ;
        RECT  13.180 3.500 13.520 3.990 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.780 1.270 14.995 3.930 ;
        RECT  14.735 1.270 14.780 3.980 ;
        RECT  14.660 1.270 14.735 1.845 ;
        RECT  14.440 3.640 14.735 3.980 ;
        RECT  14.630 1.355 14.660 1.845 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 2.940 1.840 3.305 ;
        RECT  1.300 2.690 1.635 3.305 ;
        RECT  1.295 2.690 1.300 3.030 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.775 1.185 2.435 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.290 -0.400 15.180 0.400 ;
        RECT  13.950 -0.400 14.290 0.575 ;
        RECT  12.210 -0.400 13.950 0.400 ;
        RECT  11.870 -0.400 12.210 0.575 ;
        RECT  10.690 -0.400 11.870 0.400 ;
        RECT  10.350 -0.400 10.690 1.310 ;
        RECT  6.035 -0.400 10.350 0.400 ;
        RECT  7.810 1.440 7.920 1.780 ;
        RECT  7.580 1.205 7.810 1.780 ;
        RECT  6.330 1.205 7.580 1.435 ;
        RECT  6.035 1.205 6.330 1.525 ;
        RECT  5.805 -0.400 6.035 1.525 ;
        RECT  4.190 -0.400 5.805 0.400 ;
        RECT  3.850 -0.400 4.190 0.960 ;
        RECT  1.460 -0.400 3.850 0.400 ;
        RECT  1.120 -0.400 1.460 0.575 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.100 4.640 15.180 5.440 ;
        RECT  13.760 4.465 14.100 5.440 ;
        RECT  12.760 4.640 13.760 5.440 ;
        RECT  12.420 3.620 12.760 5.440 ;
        RECT  10.740 4.640 12.420 5.440 ;
        RECT  10.400 4.070 10.740 5.440 ;
        RECT  8.400 4.640 10.400 5.440 ;
        RECT  7.460 4.070 8.400 5.440 ;
        RECT  4.330 4.640 7.460 5.440 ;
        RECT  3.990 4.465 4.330 5.440 ;
        RECT  1.605 4.640 3.990 5.440 ;
        RECT  1.195 4.390 1.605 5.440 ;
        RECT  0.000 4.640 1.195 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.420 2.495 13.950 2.835 ;
        RECT  13.100 2.495 13.420 3.140 ;
        RECT  13.080 1.250 13.100 3.140 ;
        RECT  12.800 1.250 13.080 2.795 ;
        RECT  12.770 1.250 12.800 1.550 ;
        RECT  12.430 1.210 12.770 1.550 ;
        RECT  12.455 1.825 12.560 2.110 ;
        RECT  12.225 1.825 12.455 3.295 ;
        RECT  11.925 1.825 12.225 2.055 ;
        RECT  11.480 3.065 12.225 3.295 ;
        RECT  11.695 1.595 11.925 2.055 ;
        RECT  11.390 1.595 11.695 1.825 ;
        RECT  11.140 3.065 11.480 3.940 ;
        RECT  11.390 0.970 11.450 1.310 ;
        RECT  11.110 0.970 11.390 1.825 ;
        RECT  11.325 2.140 11.380 2.480 ;
        RECT  11.040 2.140 11.325 2.505 ;
        RECT  10.540 1.595 11.110 1.825 ;
        RECT  9.915 2.275 11.040 2.505 ;
        RECT  10.255 1.595 10.540 2.045 ;
        RECT  10.200 1.705 10.255 2.045 ;
        RECT  9.915 4.000 10.030 4.340 ;
        RECT  9.905 2.275 9.915 4.340 ;
        RECT  9.685 1.285 9.905 4.340 ;
        RECT  9.675 1.285 9.685 4.285 ;
        RECT  9.280 1.285 9.675 1.515 ;
        RECT  8.940 1.230 9.280 1.570 ;
        RECT  9.150 2.500 9.260 2.840 ;
        RECT  8.920 2.500 9.150 3.840 ;
        RECT  7.525 3.610 8.920 3.840 ;
        RECT  8.535 1.830 8.915 2.170 ;
        RECT  8.305 0.675 8.535 3.375 ;
        RECT  6.605 0.675 8.305 0.905 ;
        RECT  7.760 3.145 8.305 3.375 ;
        RECT  8.005 2.020 8.060 2.410 ;
        RECT  7.720 2.020 8.005 2.415 ;
        RECT  6.645 2.180 7.720 2.415 ;
        RECT  7.295 2.705 7.525 3.840 ;
        RECT  7.165 3.610 7.295 3.840 ;
        RECT  6.935 3.610 7.165 4.365 ;
        RECT  4.790 4.135 6.935 4.365 ;
        RECT  6.415 1.825 6.645 3.385 ;
        RECT  6.265 0.635 6.605 0.975 ;
        RECT  5.575 1.825 6.415 2.055 ;
        RECT  6.110 3.155 6.415 3.385 ;
        RECT  5.880 3.155 6.110 3.820 ;
        RECT  5.760 2.440 6.100 2.780 ;
        RECT  5.770 3.480 5.880 3.820 ;
        RECT  5.355 2.495 5.760 2.725 ;
        RECT  5.370 1.655 5.575 2.055 ;
        RECT  5.355 3.480 5.410 3.820 ;
        RECT  5.345 1.140 5.370 2.055 ;
        RECT  5.125 2.435 5.355 3.820 ;
        RECT  5.140 1.140 5.345 1.885 ;
        RECT  3.825 1.655 5.140 1.885 ;
        RECT  4.990 2.435 5.125 2.665 ;
        RECT  5.070 3.480 5.125 3.820 ;
        RECT  4.600 2.115 4.990 2.665 ;
        RECT  4.755 0.770 4.870 1.110 ;
        RECT  4.560 3.945 4.790 4.365 ;
        RECT  4.525 0.770 4.755 1.420 ;
        RECT  3.675 3.945 4.560 4.175 ;
        RECT  2.825 1.190 4.525 1.420 ;
        RECT  3.485 1.655 3.825 2.080 ;
        RECT  3.465 2.935 3.675 4.355 ;
        RECT  3.445 2.395 3.465 4.355 ;
        RECT  3.235 2.395 3.445 3.165 ;
        RECT  2.155 4.125 3.445 4.355 ;
        RECT  2.905 2.395 3.235 2.625 ;
        RECT  2.775 3.480 3.110 3.840 ;
        RECT  2.675 1.995 2.905 2.625 ;
        RECT  2.485 1.160 2.825 1.500 ;
        RECT  2.545 2.965 2.775 3.840 ;
        RECT  2.335 1.995 2.675 2.225 ;
        RECT  2.370 2.965 2.545 3.195 ;
        RECT  2.100 1.270 2.485 1.500 ;
        RECT  2.140 2.460 2.370 3.195 ;
        RECT  1.925 3.745 2.155 4.355 ;
        RECT  2.100 2.460 2.140 2.690 ;
        RECT  1.870 1.270 2.100 2.690 ;
        RECT  0.600 3.745 1.925 3.975 ;
        RECT  0.545 1.100 0.850 1.440 ;
        RECT  0.545 3.520 0.600 3.975 ;
        RECT  0.315 1.100 0.545 3.975 ;
        RECT  0.260 3.520 0.315 3.975 ;
    END
END DFFRX1

MACRO DFFNSRXL
    CLASS CORE ;
    FOREIGN DFFNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.555 4.075 11.665 4.365 ;
        RECT  11.325 4.020 11.555 4.365 ;
        RECT  8.795 4.135 11.325 4.365 ;
        RECT  8.370 4.125 8.795 4.365 ;
        RECT  5.875 4.125 8.370 4.355 ;
        RECT  5.645 4.005 5.875 4.355 ;
        RECT  4.695 4.005 5.645 4.235 ;
        RECT  4.465 4.005 4.695 4.365 ;
        RECT  4.320 4.135 4.465 4.365 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 1.765 6.400 2.295 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.215 1.095 15.370 1.435 ;
        RECT  14.985 1.095 15.215 3.400 ;
        RECT  14.735 2.965 14.985 3.400 ;
        RECT  14.700 3.170 14.735 3.400 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.835 2.955 16.945 3.195 ;
        RECT  16.770 1.095 16.835 3.195 ;
        RECT  16.605 1.095 16.770 3.580 ;
        RECT  16.470 1.095 16.605 1.435 ;
        RECT  16.430 2.965 16.605 3.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.720 1.180 2.620 ;
        RECT  0.605 2.280 0.800 2.620 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.140 1.885 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.090 -0.400 17.160 0.400 ;
        RECT  15.750 -0.400 16.090 1.435 ;
        RECT  14.530 -0.400 15.750 0.400 ;
        RECT  14.190 -0.400 14.530 0.575 ;
        RECT  11.335 -0.400 14.190 0.400 ;
        RECT  10.995 -0.400 11.335 0.575 ;
        RECT  8.770 -0.400 10.995 0.400 ;
        RECT  8.430 -0.400 8.770 1.430 ;
        RECT  7.005 -0.400 8.430 0.400 ;
        RECT  6.775 -0.400 7.005 0.900 ;
        RECT  4.105 -0.400 6.775 0.400 ;
        RECT  3.765 -0.400 4.105 0.900 ;
        RECT  1.425 -0.400 3.765 0.400 ;
        RECT  1.085 -0.400 1.425 0.575 ;
        RECT  0.000 -0.400 1.085 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.950 4.640 17.160 5.440 ;
        RECT  15.610 4.090 15.950 5.440 ;
        RECT  13.450 4.640 15.610 5.440 ;
        RECT  13.110 3.395 13.450 5.440 ;
        RECT  12.285 4.640 13.110 5.440 ;
        RECT  12.055 3.395 12.285 5.440 ;
        RECT  11.370 3.395 12.055 3.625 ;
        RECT  5.415 4.640 12.055 5.440 ;
        RECT  11.010 3.310 11.370 3.625 ;
        RECT  10.785 3.395 11.010 3.625 ;
        RECT  10.555 3.395 10.785 3.845 ;
        RECT  8.845 3.615 10.555 3.845 ;
        RECT  8.615 3.515 8.845 3.845 ;
        RECT  8.375 3.515 8.615 3.745 ;
        RECT  5.075 4.465 5.415 5.440 ;
        RECT  4.090 4.640 5.075 5.440 ;
        RECT  3.750 4.465 4.090 5.440 ;
        RECT  1.100 4.640 3.750 5.440 ;
        RECT  0.760 4.465 1.100 5.440 ;
        RECT  0.000 4.640 0.760 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.860 2.145 16.330 2.375 ;
        RECT  15.630 2.145 15.860 3.860 ;
        RECT  14.430 3.630 15.630 3.860 ;
        RECT  14.430 1.170 14.540 1.510 ;
        RECT  14.200 1.170 14.430 3.860 ;
        RECT  13.830 3.395 14.200 3.735 ;
        RECT  13.645 1.825 13.875 3.165 ;
        RECT  13.485 0.980 13.735 1.320 ;
        RECT  13.025 1.825 13.645 2.055 ;
        RECT  11.890 2.935 13.645 3.165 ;
        RECT  13.395 0.630 13.485 1.320 ;
        RECT  13.255 0.630 13.395 1.265 ;
        RECT  12.155 0.630 13.255 0.860 ;
        RECT  12.795 1.090 13.025 2.055 ;
        RECT  12.595 1.090 12.795 1.320 ;
        RECT  12.070 1.855 12.300 2.230 ;
        RECT  12.135 0.630 12.155 1.235 ;
        RECT  11.925 0.630 12.135 1.290 ;
        RECT  10.945 1.855 12.070 2.085 ;
        RECT  11.795 0.950 11.925 1.290 ;
        RECT  11.660 2.615 11.890 3.165 ;
        RECT  10.835 2.615 11.660 2.845 ;
        RECT  10.715 1.250 10.945 2.085 ;
        RECT  10.295 1.250 10.715 1.480 ;
        RECT  9.425 0.720 10.585 0.950 ;
        RECT  10.065 1.250 10.295 3.360 ;
        RECT  9.995 1.250 10.065 1.535 ;
        RECT  9.655 3.130 10.065 3.360 ;
        RECT  9.765 1.195 9.995 1.535 ;
        RECT  9.425 2.485 9.750 2.715 ;
        RECT  9.195 0.720 9.425 3.280 ;
        RECT  7.915 1.660 9.195 1.890 ;
        RECT  7.940 3.050 9.195 3.280 ;
        RECT  8.635 2.125 8.865 2.605 ;
        RECT  7.455 2.125 8.635 2.355 ;
        RECT  7.470 2.590 8.225 2.820 ;
        RECT  7.710 3.050 7.940 3.800 ;
        RECT  7.685 0.670 7.915 1.890 ;
        RECT  7.475 0.670 7.685 0.900 ;
        RECT  7.240 2.590 7.470 3.840 ;
        RECT  7.225 1.135 7.455 2.355 ;
        RECT  6.335 3.610 7.240 3.840 ;
        RECT  5.745 1.135 7.225 1.365 ;
        RECT  6.755 1.635 6.985 3.375 ;
        RECT  6.570 2.805 6.755 3.375 ;
        RECT  5.595 2.805 6.570 3.035 ;
        RECT  6.105 3.535 6.335 3.840 ;
        RECT  3.325 3.535 6.105 3.765 ;
        RECT  5.515 1.135 5.745 2.575 ;
        RECT  5.505 1.135 5.515 1.435 ;
        RECT  5.310 2.345 5.515 2.575 ;
        RECT  5.165 1.095 5.505 1.435 ;
        RECT  5.080 2.345 5.310 3.305 ;
        RECT  4.550 1.695 5.225 1.925 ;
        RECT  4.065 3.075 5.080 3.305 ;
        RECT  4.320 1.600 4.550 1.925 ;
        RECT  3.600 1.600 4.320 1.830 ;
        RECT  3.835 2.065 4.065 3.305 ;
        RECT  3.595 1.300 3.600 1.830 ;
        RECT  3.365 1.290 3.595 2.965 ;
        RECT  2.935 1.290 3.365 1.530 ;
        RECT  2.835 2.735 3.365 2.965 ;
        RECT  3.095 3.535 3.325 4.280 ;
        RECT  2.350 1.770 3.120 2.110 ;
        RECT  2.355 4.050 3.095 4.280 ;
        RECT  2.650 0.900 2.935 1.530 ;
        RECT  2.605 2.735 2.835 3.820 ;
        RECT  2.595 0.900 2.650 1.240 ;
        RECT  2.350 2.930 2.355 4.280 ;
        RECT  2.125 1.505 2.350 4.280 ;
        RECT  1.785 0.675 2.170 1.040 ;
        RECT  2.120 1.505 2.125 3.480 ;
        RECT  2.075 1.505 2.120 1.790 ;
        RECT  1.995 3.020 2.120 3.480 ;
        RECT  1.735 1.450 2.075 1.790 ;
        RECT  1.520 3.020 1.995 3.250 ;
        RECT  1.480 3.835 1.805 4.390 ;
        RECT  0.465 0.810 1.785 1.040 ;
        RECT  0.480 3.835 1.480 4.065 ;
        RECT  0.480 2.925 0.535 3.265 ;
        RECT  0.250 2.925 0.480 4.065 ;
        RECT  0.235 0.810 0.465 1.770 ;
        RECT  0.195 2.925 0.250 3.265 ;
    END
END DFFNSRXL

MACRO DFFNSRX4
    CLASS CORE ;
    FOREIGN DFFNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.730 4.000 14.320 4.230 ;
        RECT  8.500 4.000 8.730 4.290 ;
        RECT  8.365 4.060 8.500 4.290 ;
        RECT  8.135 4.060 8.365 4.335 ;
        RECT  4.685 4.105 8.135 4.335 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.595 2.295 7.065 2.790 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.980 1.420 21.000 1.850 ;
        RECT  20.980 2.630 21.000 3.195 ;
        RECT  20.660 1.420 20.980 3.220 ;
        RECT  20.600 1.820 20.660 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.280 1.820 22.300 3.220 ;
        RECT  21.940 1.420 22.280 3.220 ;
        RECT  21.920 1.820 21.940 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.175 0.555 2.785 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 2.035 1.490 2.325 ;
        RECT  0.800 1.815 1.180 2.325 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.920 -0.400 23.100 0.400 ;
        RECT  22.580 -0.400 22.920 1.030 ;
        RECT  21.640 -0.400 22.580 0.400 ;
        RECT  21.300 -0.400 21.640 1.045 ;
        RECT  20.360 -0.400 21.300 0.400 ;
        RECT  20.020 -0.400 20.360 1.030 ;
        RECT  15.150 -0.400 20.020 0.400 ;
        RECT  14.810 -0.400 15.150 1.050 ;
        RECT  12.265 -0.400 14.810 0.400 ;
        RECT  11.925 -0.400 12.265 1.175 ;
        RECT  9.570 -0.400 11.925 0.400 ;
        RECT  9.340 -0.400 9.570 0.885 ;
        RECT  7.090 -0.400 9.340 0.400 ;
        RECT  6.720 -0.400 7.090 0.830 ;
        RECT  4.335 -0.400 6.720 0.400 ;
        RECT  3.995 -0.400 4.335 0.845 ;
        RECT  1.105 -0.400 3.995 0.400 ;
        RECT  0.765 -0.400 1.105 0.575 ;
        RECT  0.000 -0.400 0.765 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.920 4.640 23.100 5.440 ;
        RECT  22.580 4.035 22.920 5.440 ;
        RECT  21.640 4.640 22.580 5.440 ;
        RECT  21.300 4.035 21.640 5.440 ;
        RECT  20.360 4.640 21.300 5.440 ;
        RECT  20.020 4.035 20.360 5.440 ;
        RECT  17.610 4.640 20.020 5.440 ;
        RECT  17.270 3.640 17.610 5.440 ;
        RECT  15.550 4.640 17.270 5.440 ;
        RECT  15.320 2.920 15.550 5.440 ;
        RECT  13.345 4.640 15.320 5.440 ;
        RECT  13.005 4.465 13.345 5.440 ;
        RECT  12.190 4.640 13.005 5.440 ;
        RECT  11.850 4.465 12.190 5.440 ;
        RECT  9.525 4.640 11.850 5.440 ;
        RECT  9.185 4.465 9.525 5.440 ;
        RECT  4.410 4.640 9.185 5.440 ;
        RECT  4.070 4.465 4.410 5.440 ;
        RECT  1.085 4.640 4.070 5.440 ;
        RECT  0.745 4.465 1.085 5.440 ;
        RECT  0.000 4.640 0.745 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.605 2.210 22.835 3.740 ;
        RECT  20.295 3.510 22.605 3.740 ;
        RECT  20.065 1.670 20.295 3.740 ;
        RECT  19.545 1.670 20.065 1.900 ;
        RECT  19.260 3.400 20.065 3.740 ;
        RECT  19.065 2.160 19.750 2.500 ;
        RECT  19.315 1.440 19.545 1.900 ;
        RECT  18.900 1.375 19.065 3.015 ;
        RECT  18.835 1.375 18.900 3.610 ;
        RECT  18.050 1.375 18.835 1.605 ;
        RECT  18.670 2.785 18.835 3.610 ;
        RECT  18.485 0.675 18.715 1.030 ;
        RECT  18.560 3.085 18.670 3.610 ;
        RECT  18.370 1.860 18.600 2.260 ;
        RECT  16.330 3.085 18.560 3.315 ;
        RECT  17.330 0.675 18.485 0.905 ;
        RECT  16.110 1.860 18.370 2.090 ;
        RECT  17.680 1.205 18.050 1.605 ;
        RECT  16.705 1.375 17.680 1.605 ;
        RECT  16.990 0.675 17.330 1.050 ;
        RECT  15.875 0.675 16.990 0.905 ;
        RECT  16.475 1.140 16.705 1.605 ;
        RECT  16.265 1.140 16.475 1.370 ;
        RECT  16.220 3.085 16.330 3.600 ;
        RECT  15.990 2.455 16.220 3.600 ;
        RECT  15.825 1.860 16.110 2.155 ;
        RECT  14.830 2.455 15.990 2.685 ;
        RECT  15.765 0.675 15.875 1.290 ;
        RECT  13.680 1.925 15.825 2.155 ;
        RECT  15.645 0.675 15.765 1.605 ;
        RECT  15.535 0.950 15.645 1.605 ;
        RECT  14.375 1.375 15.535 1.605 ;
        RECT  14.755 3.535 14.985 4.410 ;
        RECT  14.600 2.455 14.830 3.305 ;
        RECT  8.195 3.535 14.755 3.765 ;
        RECT  12.755 3.075 14.600 3.305 ;
        RECT  14.145 0.970 14.375 1.605 ;
        RECT  13.450 0.875 13.680 2.155 ;
        RECT  13.285 0.875 13.450 1.105 ;
        RECT  13.290 1.925 13.450 2.155 ;
        RECT  13.060 1.925 13.290 2.845 ;
        RECT  11.520 1.405 13.220 1.635 ;
        RECT  11.055 1.925 13.060 2.155 ;
        RECT  12.525 2.385 12.755 3.305 ;
        RECT  12.320 2.385 12.525 2.615 ;
        RECT  11.290 0.675 11.520 1.635 ;
        RECT  10.280 0.675 11.290 0.905 ;
        RECT  10.890 1.755 11.055 3.135 ;
        RECT  10.825 1.220 10.890 3.135 ;
        RECT  10.660 1.220 10.825 1.985 ;
        RECT  10.515 2.905 10.825 3.135 ;
        RECT  10.280 2.300 10.590 2.530 ;
        RECT  10.050 0.675 10.280 3.195 ;
        RECT  8.660 2.965 10.050 3.195 ;
        RECT  9.530 1.530 9.760 2.325 ;
        RECT  9.110 1.530 9.530 1.760 ;
        RECT  8.880 0.935 9.110 1.760 ;
        RECT  7.735 0.935 8.880 1.165 ;
        RECT  8.560 2.565 8.660 3.195 ;
        RECT  8.560 1.400 8.650 2.000 ;
        RECT  8.430 1.400 8.560 3.195 ;
        RECT  8.420 1.400 8.430 2.795 ;
        RECT  8.330 1.765 8.420 2.795 ;
        RECT  7.965 3.085 8.195 3.765 ;
        RECT  7.605 3.085 7.965 3.315 ;
        RECT  7.605 1.530 7.780 1.760 ;
        RECT  7.505 0.935 7.735 1.295 ;
        RECT  7.680 3.605 7.735 3.835 ;
        RECT  7.450 3.605 7.680 3.840 ;
        RECT  7.375 1.530 7.605 3.315 ;
        RECT  5.695 1.065 7.505 1.295 ;
        RECT  3.830 3.610 7.450 3.840 ;
        RECT  6.170 3.085 7.375 3.315 ;
        RECT  5.940 2.280 6.170 3.315 ;
        RECT  5.465 1.065 5.695 3.375 ;
        RECT  5.400 1.065 5.465 1.435 ;
        RECT  4.130 3.145 5.465 3.375 ;
        RECT  5.005 1.755 5.235 2.240 ;
        RECT  4.755 1.755 5.005 1.985 ;
        RECT  4.525 1.565 4.755 1.985 ;
        RECT  3.600 1.565 4.525 1.795 ;
        RECT  3.900 2.330 4.130 3.375 ;
        RECT  3.600 3.610 3.830 4.410 ;
        RECT  3.370 0.785 3.600 3.080 ;
        RECT  2.835 4.180 3.600 4.410 ;
        RECT  2.840 0.785 3.370 1.015 ;
        RECT  3.300 2.850 3.370 3.080 ;
        RECT  3.070 2.850 3.300 3.825 ;
        RECT  3.080 1.750 3.135 2.090 ;
        RECT  2.795 1.750 3.080 2.100 ;
        RECT  2.605 2.905 2.835 4.410 ;
        RECT  1.975 1.755 2.795 2.100 ;
        RECT  1.975 2.905 2.605 3.135 ;
        RECT  2.265 0.725 2.460 0.955 ;
        RECT  2.055 3.735 2.370 4.170 ;
        RECT  2.035 0.725 2.265 1.045 ;
        RECT  0.520 3.820 2.055 4.050 ;
        RECT  0.545 0.815 2.035 1.045 ;
        RECT  1.745 1.425 1.975 3.360 ;
        RECT  1.565 1.425 1.745 1.655 ;
        RECT  1.525 3.020 1.745 3.360 ;
        RECT  0.315 0.815 0.545 1.635 ;
        RECT  0.290 3.210 0.520 4.050 ;
        RECT  0.205 1.295 0.315 1.635 ;
        RECT  0.180 3.210 0.290 3.550 ;
    END
END DFFNSRX4

MACRO DFFNSRX2
    CLASS CORE ;
    FOREIGN DFFNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.230 3.995 11.740 4.365 ;
        RECT  11.005 4.085 11.230 4.365 ;
        RECT  8.795 4.135 11.005 4.365 ;
        RECT  8.370 4.125 8.795 4.365 ;
        RECT  5.845 4.125 8.370 4.355 ;
        RECT  5.615 4.005 5.845 4.355 ;
        RECT  4.765 4.005 5.615 4.235 ;
        RECT  4.425 4.005 4.765 4.290 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 1.765 6.480 2.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.315 1.190 15.370 1.530 ;
        RECT  15.215 1.165 15.315 1.530 ;
        RECT  14.985 1.165 15.215 2.940 ;
        RECT  14.755 2.710 14.985 3.280 ;
        RECT  14.735 2.965 14.755 3.225 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.915 2.955 16.945 3.230 ;
        RECT  16.895 1.105 16.915 3.230 ;
        RECT  16.890 1.105 16.895 4.140 ;
        RECT  16.685 1.050 16.890 4.140 ;
        RECT  16.550 1.050 16.685 1.390 ;
        RECT  16.635 2.965 16.685 4.140 ;
        RECT  16.430 3.200 16.635 4.140 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.040 0.845 2.660 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 2.045 1.840 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.130 -0.400 17.160 0.400 ;
        RECT  15.790 -0.400 16.130 1.690 ;
        RECT  14.395 -0.400 15.790 0.400 ;
        RECT  14.055 -0.400 14.395 0.575 ;
        RECT  11.355 -0.400 14.055 0.400 ;
        RECT  11.015 -0.400 11.355 0.575 ;
        RECT  8.785 -0.400 11.015 0.400 ;
        RECT  8.445 -0.400 8.785 1.370 ;
        RECT  7.010 -0.400 8.445 0.400 ;
        RECT  6.780 -0.400 7.010 0.900 ;
        RECT  4.095 -0.400 6.780 0.400 ;
        RECT  3.755 -0.400 4.095 0.900 ;
        RECT  1.180 -0.400 3.755 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.950 4.640 17.160 5.440 ;
        RECT  15.610 4.090 15.950 5.440 ;
        RECT  13.370 4.640 15.610 5.440 ;
        RECT  13.030 3.560 13.370 5.440 ;
        RECT  12.285 4.640 13.030 5.440 ;
        RECT  12.055 3.485 12.285 5.440 ;
        RECT  10.785 3.485 12.055 3.715 ;
        RECT  5.380 4.640 12.055 5.440 ;
        RECT  10.555 3.485 10.785 3.845 ;
        RECT  8.845 3.615 10.555 3.845 ;
        RECT  8.615 3.515 8.845 3.845 ;
        RECT  8.375 3.515 8.615 3.745 ;
        RECT  5.040 4.465 5.380 5.440 ;
        RECT  4.155 4.640 5.040 5.440 ;
        RECT  3.815 4.465 4.155 5.440 ;
        RECT  1.165 4.640 3.815 5.440 ;
        RECT  0.825 4.465 1.165 5.440 ;
        RECT  0.000 4.640 0.825 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.825 2.145 16.330 2.375 ;
        RECT  15.595 2.145 15.825 3.830 ;
        RECT  14.455 3.600 15.595 3.830 ;
        RECT  14.430 3.600 14.455 3.895 ;
        RECT  14.415 1.225 14.430 3.950 ;
        RECT  14.200 1.170 14.415 3.950 ;
        RECT  14.075 1.170 14.200 1.510 ;
        RECT  14.095 3.665 14.200 3.950 ;
        RECT  13.755 3.665 14.095 4.005 ;
        RECT  13.685 1.825 13.915 3.165 ;
        RECT  12.900 1.825 13.685 2.055 ;
        RECT  11.695 2.935 13.685 3.165 ;
        RECT  13.540 0.780 13.595 1.120 ;
        RECT  13.255 0.745 13.540 1.120 ;
        RECT  12.155 0.745 13.255 0.975 ;
        RECT  12.670 1.275 12.900 2.055 ;
        RECT  12.535 1.275 12.670 1.505 ;
        RECT  12.070 1.855 12.300 2.230 ;
        RECT  11.870 0.745 12.155 1.120 ;
        RECT  10.945 1.855 12.070 2.085 ;
        RECT  11.815 0.780 11.870 1.120 ;
        RECT  11.465 2.615 11.695 3.165 ;
        RECT  10.610 2.615 11.465 2.845 ;
        RECT  10.715 1.335 10.945 2.085 ;
        RECT  10.295 1.335 10.715 1.565 ;
        RECT  9.440 0.735 10.585 0.965 ;
        RECT  10.065 1.335 10.295 3.325 ;
        RECT  9.725 1.280 10.065 1.620 ;
        RECT  9.655 3.095 10.065 3.325 ;
        RECT  9.455 2.525 9.750 2.755 ;
        RECT  9.440 1.600 9.455 2.755 ;
        RECT  9.420 0.735 9.440 2.755 ;
        RECT  9.210 0.735 9.420 3.285 ;
        RECT  7.930 1.600 9.210 1.830 ;
        RECT  9.190 2.525 9.210 3.285 ;
        RECT  7.940 3.055 9.190 3.285 ;
        RECT  8.730 2.060 8.960 2.515 ;
        RECT  7.470 2.060 8.730 2.290 ;
        RECT  7.480 2.525 8.115 2.755 ;
        RECT  7.710 3.055 7.940 3.800 ;
        RECT  7.700 0.630 7.930 1.830 ;
        RECT  7.495 0.630 7.700 0.860 ;
        RECT  7.250 2.525 7.480 3.890 ;
        RECT  7.240 1.135 7.470 2.290 ;
        RECT  6.305 3.660 7.250 3.890 ;
        RECT  5.570 1.135 7.240 1.365 ;
        RECT  6.780 1.600 7.010 3.375 ;
        RECT  6.535 2.905 6.780 3.375 ;
        RECT  5.910 2.905 6.535 3.135 ;
        RECT  6.075 3.545 6.305 3.890 ;
        RECT  3.720 3.545 6.075 3.775 ;
        RECT  5.680 2.500 5.910 3.135 ;
        RECT  5.450 1.120 5.570 1.460 ;
        RECT  5.220 1.120 5.450 3.315 ;
        RECT  3.890 3.085 5.220 3.315 ;
        RECT  4.760 1.650 4.990 2.205 ;
        RECT  3.430 1.975 4.760 2.205 ;
        RECT  3.660 2.500 3.890 3.315 ;
        RECT  3.490 3.545 3.720 3.830 ;
        RECT  2.520 3.600 3.490 3.830 ;
        RECT  3.200 1.010 3.430 2.965 ;
        RECT  2.935 1.010 3.200 1.240 ;
        RECT  2.980 2.735 3.200 2.965 ;
        RECT  2.750 2.735 2.980 3.370 ;
        RECT  2.335 1.770 2.970 2.115 ;
        RECT  2.595 0.900 2.935 1.240 ;
        RECT  2.335 3.280 2.520 3.830 ;
        RECT  2.290 1.510 2.335 3.830 ;
        RECT  2.140 1.510 2.290 3.645 ;
        RECT  2.105 1.510 2.140 3.535 ;
        RECT  1.965 1.510 2.105 1.750 ;
        RECT  1.625 3.305 2.105 3.535 ;
        RECT  1.700 0.635 2.075 1.055 ;
        RECT  1.735 3.960 2.060 4.380 ;
        RECT  1.625 1.410 1.965 1.750 ;
        RECT  0.605 3.960 1.735 4.190 ;
        RECT  0.510 0.825 1.700 1.055 ;
        RECT  0.375 3.060 0.605 4.190 ;
        RECT  0.280 0.825 0.510 1.750 ;
        RECT  0.265 3.060 0.375 3.400 ;
    END
END DFFNSRX2

MACRO DFFNSRX1
    CLASS CORE ;
    FOREIGN DFFNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.505 4.035 11.665 4.365 ;
        RECT  11.275 3.980 11.505 4.365 ;
        RECT  8.550 4.135 11.275 4.365 ;
        RECT  8.320 4.125 8.550 4.365 ;
        RECT  5.745 4.125 8.320 4.355 ;
        RECT  5.515 4.005 5.745 4.355 ;
        RECT  4.590 4.005 5.515 4.235 ;
        RECT  4.250 4.005 4.590 4.365 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.650 1.785 6.460 2.175 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.595 2.940 14.965 3.225 ;
        RECT  14.595 1.460 14.650 1.800 ;
        RECT  14.365 1.460 14.595 3.225 ;
        RECT  14.310 1.460 14.365 1.800 ;
        RECT  14.330 2.995 14.365 3.225 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.210 2.940 16.285 3.705 ;
        RECT  16.070 1.480 16.210 3.705 ;
        RECT  15.980 1.480 16.070 3.760 ;
        RECT  15.970 1.480 15.980 1.710 ;
        RECT  15.730 3.420 15.980 3.760 ;
        RECT  15.630 1.370 15.970 1.710 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.280 0.570 2.620 ;
        RECT  0.140 2.085 0.520 2.995 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.695 2.985 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.210 -0.400 16.500 0.400 ;
        RECT  14.870 -0.400 15.210 0.575 ;
        RECT  11.270 -0.400 14.870 0.400 ;
        RECT  10.930 -0.400 11.270 0.575 ;
        RECT  8.705 -0.400 10.930 0.400 ;
        RECT  8.365 -0.400 8.705 1.380 ;
        RECT  6.755 -0.400 8.365 0.400 ;
        RECT  6.525 -0.400 6.755 0.900 ;
        RECT  3.960 -0.400 6.525 0.400 ;
        RECT  3.620 -0.400 3.960 0.900 ;
        RECT  1.230 -0.400 3.620 0.400 ;
        RECT  0.890 -0.400 1.230 0.575 ;
        RECT  0.000 -0.400 0.890 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.510 4.640 16.500 5.440 ;
        RECT  15.170 4.465 15.510 5.440 ;
        RECT  13.400 4.640 15.170 5.440 ;
        RECT  13.060 3.650 13.400 5.440 ;
        RECT  12.200 4.640 13.060 5.440 ;
        RECT  11.970 3.430 12.200 5.440 ;
        RECT  10.735 3.430 11.970 3.660 ;
        RECT  5.280 4.640 11.970 5.440 ;
        RECT  10.505 3.430 10.735 3.845 ;
        RECT  8.795 3.615 10.505 3.845 ;
        RECT  8.565 3.520 8.795 3.845 ;
        RECT  8.285 3.520 8.565 3.750 ;
        RECT  4.940 4.465 5.280 5.440 ;
        RECT  4.020 4.640 4.940 5.440 ;
        RECT  3.680 4.465 4.020 5.440 ;
        RECT  1.120 4.640 3.680 5.440 ;
        RECT  0.780 4.465 1.120 5.440 ;
        RECT  0.000 4.640 0.780 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.500 2.145 15.610 2.375 ;
        RECT  15.270 2.145 15.500 3.690 ;
        RECT  13.960 3.460 15.270 3.690 ;
        RECT  13.960 0.630 14.010 2.230 ;
        RECT  13.780 0.630 13.960 3.690 ;
        RECT  13.670 0.630 13.780 0.860 ;
        RECT  13.730 2.000 13.780 3.690 ;
        RECT  13.620 2.880 13.730 3.220 ;
        RECT  12.775 2.310 13.495 2.650 ;
        RECT  13.240 1.385 13.455 1.730 ;
        RECT  13.225 0.630 13.240 1.730 ;
        RECT  13.010 0.630 13.225 1.615 ;
        RECT  12.030 0.630 13.010 0.860 ;
        RECT  12.545 1.090 12.775 3.165 ;
        RECT  12.410 1.090 12.545 1.320 ;
        RECT  11.645 2.935 12.545 3.165 ;
        RECT  11.980 1.855 12.210 2.230 ;
        RECT  11.800 0.630 12.030 1.290 ;
        RECT  10.080 1.855 11.980 2.085 ;
        RECT  11.690 0.950 11.800 1.290 ;
        RECT  11.415 2.615 11.645 3.165 ;
        RECT  10.555 2.615 11.415 2.845 ;
        RECT  10.460 0.715 10.515 0.945 ;
        RECT  10.230 0.710 10.460 0.945 ;
        RECT  9.375 0.710 10.230 0.940 ;
        RECT  9.850 1.175 10.080 3.330 ;
        RECT  9.810 1.175 9.850 2.085 ;
        RECT  9.605 3.100 9.850 3.330 ;
        RECT  9.645 1.175 9.810 1.405 ;
        RECT  9.375 2.525 9.615 2.755 ;
        RECT  9.370 0.710 9.375 2.755 ;
        RECT  9.145 0.710 9.370 3.225 ;
        RECT  7.850 1.615 9.145 1.845 ;
        RECT  9.140 2.525 9.145 3.225 ;
        RECT  7.850 2.995 9.140 3.225 ;
        RECT  8.570 2.075 8.800 2.605 ;
        RECT  7.390 2.075 8.570 2.305 ;
        RECT  7.390 2.535 8.185 2.765 ;
        RECT  7.620 0.675 7.850 1.845 ;
        RECT  7.620 2.995 7.850 3.800 ;
        RECT  7.410 0.675 7.620 0.905 ;
        RECT  7.160 1.135 7.390 2.305 ;
        RECT  7.160 2.535 7.390 3.845 ;
        RECT  5.400 1.135 7.160 1.365 ;
        RECT  6.205 3.615 7.160 3.845 ;
        RECT  6.920 2.555 6.930 2.895 ;
        RECT  6.780 1.635 6.920 2.895 ;
        RECT  6.690 1.635 6.780 3.375 ;
        RECT  6.495 2.555 6.690 3.375 ;
        RECT  6.440 2.905 6.495 3.375 ;
        RECT  5.775 2.905 6.440 3.135 ;
        RECT  5.975 3.515 6.205 3.845 ;
        RECT  3.315 3.515 5.975 3.745 ;
        RECT  5.545 2.540 5.775 3.135 ;
        RECT  5.315 1.120 5.400 1.460 ;
        RECT  5.085 1.120 5.315 3.135 ;
        RECT  5.060 1.120 5.085 1.460 ;
        RECT  4.820 2.905 5.085 3.135 ;
        RECT  4.625 1.840 4.855 2.205 ;
        RECT  3.755 2.905 4.820 3.260 ;
        RECT  3.295 1.975 4.625 2.205 ;
        RECT  3.525 2.510 3.755 3.260 ;
        RECT  3.085 3.515 3.315 4.410 ;
        RECT  3.065 0.955 3.295 2.965 ;
        RECT  2.385 4.180 3.085 4.410 ;
        RECT  2.730 0.955 3.065 1.240 ;
        RECT  2.845 2.735 3.065 2.965 ;
        RECT  2.615 2.735 2.845 3.525 ;
        RECT  2.385 1.770 2.835 2.110 ;
        RECT  2.390 0.900 2.730 1.240 ;
        RECT  2.155 1.485 2.385 4.410 ;
        RECT  1.920 1.485 2.155 1.720 ;
        RECT  1.540 3.250 2.155 3.535 ;
        RECT  1.690 0.695 1.930 0.925 ;
        RECT  1.600 4.005 1.925 4.380 ;
        RECT  1.580 1.380 1.920 1.720 ;
        RECT  1.460 0.695 1.690 1.040 ;
        RECT  0.520 4.005 1.600 4.235 ;
        RECT  0.465 0.810 1.460 1.040 ;
        RECT  0.290 3.400 0.520 4.235 ;
        RECT  0.235 0.810 0.465 1.720 ;
        RECT  0.180 3.400 0.290 3.740 ;
    END
END DFFNSRX1

MACRO DFFNSXL
    CLASS CORE ;
    FOREIGN DFFNSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 3.770 10.675 4.340 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.655 0.865 12.885 3.755 ;
        RECT  12.255 0.865 12.655 1.095 ;
        RECT  12.395 3.500 12.655 3.755 ;
        RECT  12.325 3.525 12.395 3.755 ;
        RECT  12.095 3.525 12.325 3.850 ;
        RECT  12.025 0.745 12.255 1.095 ;
        RECT  12.070 3.620 12.095 3.850 ;
        RECT  11.840 3.620 12.070 4.195 ;
        RECT  11.500 0.745 12.025 0.975 ;
        RECT  11.730 3.855 11.840 4.195 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.420 1.210 13.660 3.250 ;
        RECT  13.340 1.210 13.420 3.435 ;
        RECT  13.185 1.210 13.340 1.590 ;
        RECT  13.165 2.845 13.340 3.435 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.370 1.840 2.095 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.685 2.280 1.180 2.700 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.870 -0.400 13.860 0.400 ;
        RECT  12.530 -0.400 12.870 0.575 ;
        RECT  11.100 -0.400 12.530 0.400 ;
        RECT  10.760 -0.400 11.100 1.030 ;
        RECT  9.040 -0.400 10.760 0.400 ;
        RECT  8.700 -0.400 9.040 0.575 ;
        RECT  6.470 -0.400 8.700 0.400 ;
        RECT  6.240 -0.400 6.470 1.135 ;
        RECT  4.160 -0.400 6.240 0.400 ;
        RECT  3.820 -0.400 4.160 1.065 ;
        RECT  1.275 -0.400 3.820 0.400 ;
        RECT  0.935 -0.400 1.275 0.575 ;
        RECT  0.000 -0.400 0.935 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.930 4.640 13.860 5.440 ;
        RECT  12.495 4.465 12.930 5.440 ;
        RECT  11.235 4.640 12.495 5.440 ;
        RECT  11.005 3.265 11.235 5.440 ;
        RECT  9.680 4.640 11.005 5.440 ;
        RECT  9.340 4.140 9.680 5.440 ;
        RECT  7.090 4.640 9.340 5.440 ;
        RECT  6.860 3.765 7.090 5.440 ;
        RECT  5.695 4.640 6.860 5.440 ;
        RECT  5.355 4.110 5.695 5.440 ;
        RECT  4.405 4.640 5.355 5.440 ;
        RECT  4.065 4.465 4.405 5.440 ;
        RECT  1.470 4.640 4.065 5.440 ;
        RECT  1.130 4.465 1.470 5.440 ;
        RECT  0.000 4.640 1.130 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.155 1.600 12.185 2.375 ;
        RECT  11.955 1.600 12.155 3.190 ;
        RECT  11.880 1.600 11.955 1.830 ;
        RECT  11.925 2.075 11.955 3.190 ;
        RECT  11.710 2.960 11.925 3.190 ;
        RECT  11.540 1.490 11.880 1.830 ;
        RECT  11.110 2.140 11.450 2.480 ;
        RECT  10.515 2.195 11.110 2.425 ;
        RECT  10.490 1.620 10.515 3.375 ;
        RECT  10.285 1.620 10.490 3.430 ;
        RECT  9.740 1.620 10.285 1.850 ;
        RECT  10.150 3.090 10.285 3.430 ;
        RECT  8.500 2.435 10.030 2.665 ;
        RECT  9.400 1.190 9.740 1.850 ;
        RECT  9.210 1.620 9.400 1.850 ;
        RECT  8.870 1.620 9.210 1.960 ;
        RECT  8.465 1.545 8.500 3.835 ;
        RECT  8.270 1.545 8.465 3.890 ;
        RECT  7.215 0.675 8.290 0.905 ;
        RECT  7.825 1.545 8.270 1.775 ;
        RECT  8.125 3.550 8.270 3.890 ;
        RECT  7.215 2.515 8.040 2.915 ;
        RECT  7.595 1.190 7.825 1.775 ;
        RECT  6.985 0.675 7.215 2.915 ;
        RECT  6.010 1.370 6.985 1.600 ;
        RECT  6.445 2.685 6.985 2.915 ;
        RECT  5.795 1.855 6.755 2.085 ;
        RECT  6.215 2.685 6.445 3.405 ;
        RECT  5.945 3.650 6.175 4.040 ;
        RECT  5.780 0.695 6.010 1.600 ;
        RECT  3.610 3.650 5.945 3.880 ;
        RECT  5.565 1.855 5.795 3.415 ;
        RECT  4.710 0.630 5.780 0.925 ;
        RECT  5.550 1.855 5.565 2.085 ;
        RECT  4.465 3.185 5.565 3.415 ;
        RECT  5.320 1.450 5.550 2.085 ;
        RECT  5.095 2.355 5.325 2.740 ;
        RECT  4.985 2.355 5.095 2.585 ;
        RECT  4.755 1.320 4.985 2.585 ;
        RECT  3.575 1.320 4.755 1.550 ;
        RECT  4.655 0.630 4.710 0.860 ;
        RECT  4.235 2.035 4.465 3.415 ;
        RECT  3.755 2.035 4.235 2.265 ;
        RECT  3.380 2.570 3.610 4.205 ;
        RECT  3.345 1.130 3.575 1.550 ;
        RECT  3.305 2.570 3.380 2.800 ;
        RECT  1.960 3.975 3.380 4.205 ;
        RECT  2.795 1.130 3.345 1.360 ;
        RECT  3.105 1.885 3.305 2.800 ;
        RECT  2.895 3.035 3.125 3.520 ;
        RECT  3.075 1.600 3.105 2.800 ;
        RECT  2.820 1.600 3.075 2.115 ;
        RECT  2.840 3.035 2.895 3.265 ;
        RECT  2.610 2.595 2.840 3.265 ;
        RECT  2.505 0.870 2.795 1.360 ;
        RECT  2.505 2.595 2.610 2.825 ;
        RECT  2.455 0.870 2.505 2.825 ;
        RECT  2.275 1.130 2.455 2.825 ;
        RECT  1.730 3.945 1.960 4.205 ;
        RECT  0.395 3.945 1.730 4.175 ;
        RECT  0.395 1.195 0.540 1.535 ;
        RECT  0.395 3.295 0.520 3.635 ;
        RECT  0.200 1.195 0.395 4.175 ;
        RECT  0.165 1.225 0.200 4.175 ;
    END
END DFFNSXL

MACRO DFFNSX4
    CLASS CORE ;
    FOREIGN DFFNSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.470 4.010 5.090 4.390 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.020 2.875 17.035 3.215 ;
        RECT  16.800 1.200 17.020 3.215 ;
        RECT  16.695 0.715 16.800 3.215 ;
        RECT  16.640 0.715 16.695 2.660 ;
        RECT  16.460 0.715 16.640 1.655 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.340 0.955 18.350 2.700 ;
        RECT  18.240 0.955 18.340 3.220 ;
        RECT  17.960 0.760 18.240 3.220 ;
        RECT  17.955 0.760 17.960 3.160 ;
        RECT  17.900 0.760 17.955 1.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.590 1.445 1.930 2.090 ;
        RECT  1.535 1.835 1.590 2.075 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 2.055 1.170 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.960 -0.400 19.140 0.400 ;
        RECT  18.620 -0.400 18.960 1.565 ;
        RECT  17.520 -0.400 18.620 0.400 ;
        RECT  17.180 -0.400 17.520 0.960 ;
        RECT  16.040 -0.400 17.180 0.400 ;
        RECT  15.700 -0.400 16.040 0.915 ;
        RECT  14.780 -0.400 15.700 0.400 ;
        RECT  14.440 -0.400 14.780 1.190 ;
        RECT  12.175 -0.400 14.440 0.400 ;
        RECT  11.835 -0.400 12.175 0.575 ;
        RECT  10.100 -0.400 11.835 0.400 ;
        RECT  9.760 -0.400 10.100 0.575 ;
        RECT  7.420 -0.400 9.760 0.400 ;
        RECT  7.080 -0.400 7.420 1.080 ;
        RECT  4.375 -0.400 7.080 0.400 ;
        RECT  4.035 -0.400 4.375 1.225 ;
        RECT  1.395 -0.400 4.035 0.400 ;
        RECT  1.055 -0.400 1.395 0.575 ;
        RECT  0.000 -0.400 1.055 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.955 4.640 19.140 5.440 ;
        RECT  18.615 4.055 18.955 5.440 ;
        RECT  17.675 4.640 18.615 5.440 ;
        RECT  17.335 4.015 17.675 5.440 ;
        RECT  16.395 4.640 17.335 5.440 ;
        RECT  16.055 4.055 16.395 5.440 ;
        RECT  14.970 4.640 16.055 5.440 ;
        RECT  14.630 3.520 14.970 5.440 ;
        RECT  13.530 4.640 14.630 5.440 ;
        RECT  13.190 3.520 13.530 5.440 ;
        RECT  12.050 4.640 13.190 5.440 ;
        RECT  11.710 4.015 12.050 5.440 ;
        RECT  9.980 4.640 11.710 5.440 ;
        RECT  9.640 3.380 9.980 5.440 ;
        RECT  7.380 4.640 9.640 5.440 ;
        RECT  7.040 3.330 7.380 5.440 ;
        RECT  5.720 4.640 7.040 5.440 ;
        RECT  5.380 4.195 5.720 5.440 ;
        RECT  4.175 4.640 5.380 5.440 ;
        RECT  3.945 4.150 4.175 5.440 ;
        RECT  1.390 4.640 3.945 5.440 ;
        RECT  1.050 4.465 1.390 5.440 ;
        RECT  0.000 4.640 1.050 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.645 2.060 18.875 3.725 ;
        RECT  16.115 3.495 18.645 3.725 ;
        RECT  15.885 1.620 16.115 3.725 ;
        RECT  15.500 1.620 15.885 1.850 ;
        RECT  15.690 3.055 15.885 3.725 ;
        RECT  15.350 3.055 15.690 3.865 ;
        RECT  15.215 1.280 15.500 1.850 ;
        RECT  14.250 2.080 15.460 2.420 ;
        RECT  15.160 1.280 15.215 1.620 ;
        RECT  14.195 2.080 14.250 3.340 ;
        RECT  14.020 1.505 14.195 3.340 ;
        RECT  13.965 1.505 14.020 2.310 ;
        RECT  13.910 2.975 14.020 3.340 ;
        RECT  13.590 1.505 13.965 1.735 ;
        RECT  12.810 2.975 13.910 3.205 ;
        RECT  13.280 2.130 13.620 2.470 ;
        RECT  13.525 1.295 13.590 1.735 ;
        RECT  13.360 1.055 13.525 1.735 ;
        RECT  13.160 1.055 13.360 1.580 ;
        RECT  10.855 2.185 13.280 2.415 ;
        RECT  11.435 1.055 13.160 1.285 ;
        RECT  12.700 2.975 12.810 3.340 ;
        RECT  12.470 2.975 12.700 3.725 ;
        RECT  11.460 3.495 12.470 3.725 ;
        RECT  11.230 3.495 11.460 4.040 ;
        RECT  9.405 0.865 10.975 1.095 ;
        RECT  10.630 1.385 10.855 3.085 ;
        RECT  10.625 1.385 10.630 3.260 ;
        RECT  10.355 1.385 10.625 1.770 ;
        RECT  10.400 2.855 10.625 3.260 ;
        RECT  8.660 2.915 10.400 3.145 ;
        RECT  10.080 2.275 10.390 2.505 ;
        RECT  8.940 1.385 10.355 1.615 ;
        RECT  9.850 2.175 10.080 2.505 ;
        RECT  9.505 2.175 9.850 2.405 ;
        RECT  9.275 1.925 9.505 2.405 ;
        RECT  9.175 0.675 9.405 1.095 ;
        RECT  8.740 1.925 9.275 2.155 ;
        RECT  8.100 0.675 9.175 0.905 ;
        RECT  8.710 1.195 8.940 1.615 ;
        RECT  8.400 1.195 8.710 1.425 ;
        RECT  8.375 2.915 8.660 3.440 ;
        RECT  8.015 2.310 8.410 2.650 ;
        RECT  8.320 3.100 8.375 3.440 ;
        RECT  8.015 0.675 8.100 1.625 ;
        RECT  7.870 0.675 8.015 3.100 ;
        RECT  7.785 1.395 7.870 3.100 ;
        RECT  6.620 1.395 7.785 1.645 ;
        RECT  6.705 2.870 7.785 3.100 ;
        RECT  6.215 2.235 7.495 2.635 ;
        RECT  6.475 2.870 6.705 3.265 ;
        RECT  6.335 0.675 6.620 1.645 ;
        RECT  6.105 3.035 6.475 3.265 ;
        RECT  6.115 3.520 6.345 4.100 ;
        RECT  6.280 0.675 6.335 1.600 ;
        RECT  6.180 0.675 6.280 1.040 ;
        RECT  5.815 2.230 6.215 2.635 ;
        RECT  3.515 3.520 6.115 3.750 ;
        RECT  5.710 1.715 5.815 3.265 ;
        RECT  5.585 1.015 5.710 3.265 ;
        RECT  5.480 1.015 5.585 1.945 ;
        RECT  4.090 3.035 5.585 3.265 ;
        RECT  5.315 1.015 5.480 1.245 ;
        RECT  5.005 2.455 5.290 2.685 ;
        RECT  4.775 1.495 5.005 2.685 ;
        RECT  3.015 1.495 4.775 1.725 ;
        RECT  3.860 2.010 4.090 3.265 ;
        RECT  3.285 2.075 3.515 4.345 ;
        RECT  3.065 2.075 3.285 2.305 ;
        RECT  1.885 4.115 3.285 4.345 ;
        RECT  2.835 3.000 3.050 3.710 ;
        RECT  2.905 1.000 3.015 1.725 ;
        RECT  2.835 1.000 2.905 1.840 ;
        RECT  2.820 1.000 2.835 3.710 ;
        RECT  2.675 1.000 2.820 3.230 ;
        RECT  2.605 1.610 2.675 3.230 ;
        RECT  1.655 3.875 1.885 4.345 ;
        RECT  0.465 3.875 1.655 4.105 ;
        RECT  0.465 1.270 0.520 1.610 ;
        RECT  0.465 2.960 0.520 3.300 ;
        RECT  0.235 1.270 0.465 4.105 ;
        RECT  0.180 1.270 0.235 1.610 ;
        RECT  0.180 2.960 0.235 3.300 ;
    END
END DFFNSX4

MACRO DFFNSX2
    CLASS CORE ;
    FOREIGN DFFNSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.760 3.950 10.405 4.405 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.145 0.835 12.325 2.920 ;
        RECT  12.130 0.690 12.145 2.920 ;
        RECT  12.095 0.690 12.130 3.110 ;
        RECT  11.915 0.690 12.095 1.065 ;
        RECT  12.020 2.635 12.095 3.110 ;
        RECT  11.900 2.690 12.020 3.110 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 1.845 13.720 3.130 ;
        RECT  13.640 0.955 13.645 3.130 ;
        RECT  13.575 0.755 13.640 3.130 ;
        RECT  13.490 0.755 13.575 4.240 ;
        RECT  13.415 0.755 13.490 2.075 ;
        RECT  13.345 2.900 13.490 4.240 ;
        RECT  13.300 0.755 13.415 1.565 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.380 1.840 1.970 ;
        RECT  1.535 1.380 1.765 2.075 ;
        RECT  1.320 1.380 1.535 1.970 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.660 2.320 1.180 2.840 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.920 -0.400 13.860 0.400 ;
        RECT  12.580 -0.400 12.920 1.475 ;
        RECT  11.060 -0.400 12.580 0.400 ;
        RECT  10.720 -0.400 11.060 0.575 ;
        RECT  9.040 -0.400 10.720 0.400 ;
        RECT  8.700 -0.400 9.040 0.575 ;
        RECT  6.470 -0.400 8.700 0.400 ;
        RECT  6.240 -0.400 6.470 1.135 ;
        RECT  4.160 -0.400 6.240 0.400 ;
        RECT  3.820 -0.400 4.160 1.065 ;
        RECT  1.400 -0.400 3.820 0.400 ;
        RECT  1.060 -0.400 1.400 0.575 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.910 4.640 13.860 5.440 ;
        RECT  12.570 3.925 12.910 5.440 ;
        RECT  10.895 4.640 12.570 5.440 ;
        RECT  10.865 3.505 10.895 5.440 ;
        RECT  10.665 3.340 10.865 5.440 ;
        RECT  10.635 3.340 10.665 3.735 ;
        RECT  9.440 4.640 10.665 5.440 ;
        RECT  9.100 4.140 9.440 5.440 ;
        RECT  6.945 4.640 9.100 5.440 ;
        RECT  6.715 3.770 6.945 5.440 ;
        RECT  5.695 4.640 6.715 5.440 ;
        RECT  5.355 4.095 5.695 5.440 ;
        RECT  4.405 4.640 5.355 5.440 ;
        RECT  4.065 4.465 4.405 5.440 ;
        RECT  1.440 4.640 4.065 5.440 ;
        RECT  1.100 4.465 1.440 5.440 ;
        RECT  0.000 4.640 1.100 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.110 2.240 13.150 2.620 ;
        RECT  12.920 2.240 13.110 3.585 ;
        RECT  12.880 2.295 12.920 3.585 ;
        RECT  11.615 3.355 12.880 3.585 ;
        RECT  11.615 1.435 11.655 1.775 ;
        RECT  11.590 1.435 11.615 3.585 ;
        RECT  11.385 1.435 11.590 3.830 ;
        RECT  11.315 1.435 11.385 1.775 ;
        RECT  11.360 3.355 11.385 3.830 ;
        RECT  10.380 2.120 11.155 2.505 ;
        RECT  10.200 1.620 10.380 3.125 ;
        RECT  10.150 1.620 10.200 3.635 ;
        RECT  9.740 1.620 10.150 1.850 ;
        RECT  9.860 2.825 10.150 3.635 ;
        RECT  8.315 2.195 9.920 2.425 ;
        RECT  9.400 1.160 9.740 1.850 ;
        RECT  9.010 1.620 9.400 1.850 ;
        RECT  8.670 1.620 9.010 1.960 ;
        RECT  8.280 1.545 8.315 3.835 ;
        RECT  7.215 0.675 8.290 0.905 ;
        RECT  8.085 1.545 8.280 3.890 ;
        RECT  7.825 1.545 8.085 1.775 ;
        RECT  7.940 3.550 8.085 3.890 ;
        RECT  7.215 2.515 7.855 2.915 ;
        RECT  7.595 1.190 7.825 1.775 ;
        RECT  6.985 0.675 7.215 2.915 ;
        RECT  6.010 1.370 6.985 1.600 ;
        RECT  6.405 2.685 6.985 2.915 ;
        RECT  6.515 1.885 6.745 2.295 ;
        RECT  5.795 1.885 6.515 2.115 ;
        RECT  6.175 2.685 6.405 3.405 ;
        RECT  5.945 3.635 6.175 4.040 ;
        RECT  5.780 0.695 6.010 1.600 ;
        RECT  3.610 3.635 5.945 3.865 ;
        RECT  5.565 1.885 5.795 3.370 ;
        RECT  5.080 0.695 5.780 0.925 ;
        RECT  5.550 1.885 5.565 2.115 ;
        RECT  4.465 3.140 5.565 3.370 ;
        RECT  5.320 1.450 5.550 2.115 ;
        RECT  5.095 2.370 5.325 2.790 ;
        RECT  4.985 2.370 5.095 2.600 ;
        RECT  4.655 0.630 5.080 0.925 ;
        RECT  4.755 1.295 4.985 2.600 ;
        RECT  2.795 1.295 4.755 1.525 ;
        RECT  4.235 2.035 4.465 3.370 ;
        RECT  3.755 2.035 4.235 2.265 ;
        RECT  3.380 2.570 3.610 4.085 ;
        RECT  3.305 2.570 3.380 2.800 ;
        RECT  0.540 3.855 3.380 4.085 ;
        RECT  3.075 1.805 3.305 2.800 ;
        RECT  2.895 3.035 3.125 3.520 ;
        RECT  2.820 1.805 3.075 2.035 ;
        RECT  2.840 3.035 2.895 3.265 ;
        RECT  2.610 2.595 2.840 3.265 ;
        RECT  2.505 0.860 2.795 1.525 ;
        RECT  2.505 2.595 2.610 2.825 ;
        RECT  2.455 0.860 2.505 2.825 ;
        RECT  2.275 1.295 2.455 2.825 ;
        RECT  0.430 0.815 0.540 1.155 ;
        RECT  0.430 3.400 0.540 4.085 ;
        RECT  0.200 0.815 0.430 4.085 ;
    END
END DFFNSX2

MACRO DFFNSX1
    CLASS CORE ;
    FOREIGN DFFNSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 3.770 10.675 4.340 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.615 0.865 12.845 3.755 ;
        RECT  12.215 0.865 12.615 1.095 ;
        RECT  12.395 3.500 12.615 3.755 ;
        RECT  12.325 3.525 12.395 3.755 ;
        RECT  12.095 3.525 12.325 3.850 ;
        RECT  11.985 0.790 12.215 1.095 ;
        RECT  12.070 3.620 12.095 3.850 ;
        RECT  11.840 3.620 12.070 4.195 ;
        RECT  11.460 0.790 11.985 1.020 ;
        RECT  11.730 3.855 11.840 4.195 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.415 1.210 13.660 3.250 ;
        RECT  13.340 1.210 13.415 3.670 ;
        RECT  13.185 1.210 13.340 1.590 ;
        RECT  13.185 2.845 13.340 3.670 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.375 1.840 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.685 2.280 1.180 2.700 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.870 -0.400 13.860 0.400 ;
        RECT  12.530 -0.400 12.870 0.575 ;
        RECT  11.060 -0.400 12.530 0.400 ;
        RECT  10.720 -0.400 11.060 1.010 ;
        RECT  9.040 -0.400 10.720 0.400 ;
        RECT  8.700 -0.400 9.040 0.575 ;
        RECT  6.460 -0.400 8.700 0.400 ;
        RECT  6.230 -0.400 6.460 1.135 ;
        RECT  4.160 -0.400 6.230 0.400 ;
        RECT  3.820 -0.400 4.160 1.065 ;
        RECT  1.240 -0.400 3.820 0.400 ;
        RECT  0.900 -0.400 1.240 0.575 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.930 4.640 13.860 5.440 ;
        RECT  12.495 4.465 12.930 5.440 ;
        RECT  11.235 4.640 12.495 5.440 ;
        RECT  11.005 3.030 11.235 5.440 ;
        RECT  9.680 4.640 11.005 5.440 ;
        RECT  9.340 4.140 9.680 5.440 ;
        RECT  7.090 4.640 9.340 5.440 ;
        RECT  6.860 3.765 7.090 5.440 ;
        RECT  5.695 4.640 6.860 5.440 ;
        RECT  5.355 4.095 5.695 5.440 ;
        RECT  4.405 4.640 5.355 5.440 ;
        RECT  4.065 4.465 4.405 5.440 ;
        RECT  1.560 4.640 4.065 5.440 ;
        RECT  1.220 4.465 1.560 5.440 ;
        RECT  0.000 4.640 1.220 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.155 2.020 12.185 2.375 ;
        RECT  11.925 1.600 12.155 3.095 ;
        RECT  11.840 1.600 11.925 1.830 ;
        RECT  11.710 2.865 11.925 3.095 ;
        RECT  11.500 1.490 11.840 1.830 ;
        RECT  11.110 2.140 11.450 2.480 ;
        RECT  10.515 2.195 11.110 2.425 ;
        RECT  10.490 1.620 10.515 3.345 ;
        RECT  10.285 1.620 10.490 3.400 ;
        RECT  9.740 1.620 10.285 1.850 ;
        RECT  10.150 3.060 10.285 3.400 ;
        RECT  8.500 2.435 10.030 2.665 ;
        RECT  9.400 1.190 9.740 1.850 ;
        RECT  9.210 1.620 9.400 1.850 ;
        RECT  8.870 1.620 9.210 1.960 ;
        RECT  8.465 1.545 8.500 3.835 ;
        RECT  8.270 1.545 8.465 3.890 ;
        RECT  7.215 0.675 8.290 0.905 ;
        RECT  7.825 1.545 8.270 1.775 ;
        RECT  8.125 3.550 8.270 3.890 ;
        RECT  7.215 2.515 8.040 2.915 ;
        RECT  7.595 1.190 7.825 1.775 ;
        RECT  6.985 0.675 7.215 2.915 ;
        RECT  6.000 1.370 6.985 1.600 ;
        RECT  6.445 2.685 6.985 2.915 ;
        RECT  5.795 1.835 6.745 2.065 ;
        RECT  6.215 2.685 6.445 3.405 ;
        RECT  5.945 3.635 6.175 4.040 ;
        RECT  5.780 0.695 6.000 1.600 ;
        RECT  3.610 3.635 5.945 3.865 ;
        RECT  5.565 1.835 5.795 3.370 ;
        RECT  5.770 0.675 5.780 1.600 ;
        RECT  4.710 0.675 5.770 0.925 ;
        RECT  5.540 1.835 5.565 2.065 ;
        RECT  4.465 3.140 5.565 3.370 ;
        RECT  5.310 1.420 5.540 2.065 ;
        RECT  5.095 2.355 5.325 2.740 ;
        RECT  4.985 2.355 5.095 2.585 ;
        RECT  4.755 1.295 4.985 2.585 ;
        RECT  2.795 1.295 4.755 1.525 ;
        RECT  4.655 0.675 4.710 0.905 ;
        RECT  4.235 2.005 4.465 3.370 ;
        RECT  3.705 2.005 4.235 2.235 ;
        RECT  3.380 2.570 3.610 4.085 ;
        RECT  3.305 2.570 3.380 2.800 ;
        RECT  1.575 3.855 3.380 4.085 ;
        RECT  3.075 1.805 3.305 2.800 ;
        RECT  2.895 3.035 3.125 3.520 ;
        RECT  2.820 1.805 3.075 2.035 ;
        RECT  2.840 3.035 2.895 3.265 ;
        RECT  2.610 2.595 2.840 3.265 ;
        RECT  2.505 0.860 2.795 1.525 ;
        RECT  2.505 2.595 2.610 2.825 ;
        RECT  2.455 0.860 2.505 2.825 ;
        RECT  2.275 1.295 2.455 2.825 ;
        RECT  1.345 3.855 1.575 4.175 ;
        RECT  0.395 3.945 1.345 4.175 ;
        RECT  0.395 1.195 0.540 1.535 ;
        RECT  0.395 3.360 0.520 3.700 ;
        RECT  0.200 1.195 0.395 4.175 ;
        RECT  0.165 1.225 0.200 4.175 ;
    END
END DFFNSX1

MACRO DFFNRXL
    CLASS CORE ;
    FOREIGN DFFNRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.590 2.900 4.930 3.240 ;
        RECT  4.480 2.900 4.590 3.185 ;
        RECT  4.250 2.360 4.480 3.185 ;
        RECT  4.120 2.360 4.250 2.680 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.125 0.865 14.355 4.035 ;
        RECT  13.770 0.865 14.125 1.095 ;
        RECT  13.975 3.500 14.125 4.035 ;
        RECT  13.850 3.805 13.975 4.035 ;
        RECT  13.510 3.805 13.850 4.230 ;
        RECT  13.430 0.635 13.770 1.095 ;
        RECT  13.470 3.805 13.510 4.175 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.495 3.620 15.580 3.960 ;
        RECT  15.265 1.890 15.495 3.960 ;
        RECT  15.180 1.890 15.265 2.120 ;
        RECT  15.240 3.620 15.265 3.960 ;
        RECT  14.660 1.190 15.180 2.120 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.525 1.575 1.915 2.105 ;
        RECT  1.455 1.715 1.525 2.080 ;
        RECT  1.400 1.740 1.455 2.080 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 2.635 1.230 3.220 ;
        RECT  0.910 1.885 1.020 2.405 ;
        RECT  0.680 1.885 0.910 3.220 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.500 -0.400 15.840 0.400 ;
        RECT  14.160 -0.400 14.500 0.575 ;
        RECT  12.890 -0.400 14.160 0.400 ;
        RECT  12.550 -0.400 12.890 0.950 ;
        RECT  11.130 -0.400 12.550 0.400 ;
        RECT  10.790 -0.400 11.130 1.110 ;
        RECT  6.365 -0.400 10.790 0.400 ;
        RECT  7.895 1.205 8.235 1.760 ;
        RECT  6.660 1.205 7.895 1.435 ;
        RECT  6.365 1.205 6.660 1.580 ;
        RECT  6.320 -0.400 6.365 1.580 ;
        RECT  6.135 -0.400 6.320 1.525 ;
        RECT  4.350 -0.400 6.135 0.400 ;
        RECT  4.010 -0.400 4.350 0.960 ;
        RECT  1.350 -0.400 4.010 0.400 ;
        RECT  1.010 -0.400 1.350 0.575 ;
        RECT  0.000 -0.400 1.010 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.810 4.640 15.840 5.440 ;
        RECT  14.470 4.465 14.810 5.440 ;
        RECT  13.090 4.640 14.470 5.440 ;
        RECT  12.750 4.110 13.090 5.440 ;
        RECT  11.065 4.640 12.750 5.440 ;
        RECT  10.725 4.080 11.065 5.440 ;
        RECT  8.730 4.640 10.725 5.440 ;
        RECT  7.790 4.080 8.730 5.440 ;
        RECT  4.660 4.640 7.790 5.440 ;
        RECT  4.320 4.465 4.660 5.440 ;
        RECT  1.650 4.640 4.320 5.440 ;
        RECT  1.310 4.080 1.650 5.440 ;
        RECT  0.000 4.640 1.310 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.740 1.380 13.850 3.160 ;
        RECT  13.510 1.380 13.740 3.350 ;
        RECT  13.330 1.380 13.510 1.850 ;
        RECT  13.400 2.820 13.510 3.350 ;
        RECT  12.985 1.880 13.030 2.220 ;
        RECT  12.975 1.865 12.985 2.220 ;
        RECT  12.475 1.865 12.975 2.245 ;
        RECT  12.245 1.865 12.475 3.850 ;
        RECT  12.035 1.865 12.245 2.095 ;
        RECT  11.770 3.620 12.245 3.850 ;
        RECT  11.805 0.915 12.035 2.095 ;
        RECT  11.670 3.005 12.010 3.390 ;
        RECT  11.645 0.915 11.805 1.825 ;
        RECT  11.430 3.620 11.770 3.960 ;
        RECT  10.535 3.160 11.670 3.390 ;
        RECT  11.235 1.595 11.645 1.825 ;
        RECT  11.235 2.240 11.290 2.580 ;
        RECT  11.005 1.595 11.235 2.580 ;
        RECT  10.950 2.240 11.005 2.580 ;
        RECT  10.355 1.425 10.535 3.405 ;
        RECT  10.355 4.000 10.360 4.340 ;
        RECT  10.305 1.425 10.355 4.340 ;
        RECT  9.590 1.425 10.305 1.655 ;
        RECT  10.125 3.160 10.305 4.340 ;
        RECT  10.020 4.000 10.125 4.340 ;
        RECT  9.615 2.390 9.955 2.730 ;
        RECT  9.530 0.630 9.870 0.970 ;
        RECT  8.935 2.445 9.615 2.675 ;
        RECT  9.305 1.290 9.590 1.655 ;
        RECT  8.935 0.685 9.530 0.915 ;
        RECT  9.250 1.290 9.305 1.630 ;
        RECT  8.705 0.675 8.935 3.465 ;
        RECT  7.315 0.675 8.705 0.915 ;
        RECT  8.150 3.075 8.705 3.465 ;
        RECT  6.975 2.140 8.390 2.480 ;
        RECT  7.855 2.810 7.910 3.150 ;
        RECT  7.625 2.810 7.855 3.825 ;
        RECT  7.570 2.810 7.625 3.150 ;
        RECT  7.495 3.595 7.625 3.825 ;
        RECT  7.265 3.595 7.495 4.365 ;
        RECT  7.030 0.675 7.315 0.905 ;
        RECT  5.125 4.135 7.265 4.365 ;
        RECT  6.690 0.635 7.030 0.975 ;
        RECT  6.745 1.825 6.975 3.690 ;
        RECT  5.710 1.825 6.745 2.055 ;
        RECT  6.440 3.460 6.745 3.690 ;
        RECT  6.100 3.460 6.440 3.800 ;
        RECT  6.090 2.440 6.430 2.780 ;
        RECT  5.485 2.495 6.090 2.725 ;
        RECT  5.710 1.100 5.720 1.440 ;
        RECT  5.480 1.100 5.710 2.055 ;
        RECT  5.485 3.485 5.705 3.870 ;
        RECT  5.365 2.435 5.485 3.870 ;
        RECT  5.380 1.100 5.480 1.885 ;
        RECT  3.900 1.655 5.380 1.885 ;
        RECT  5.255 2.435 5.365 3.715 ;
        RECT  5.250 2.435 5.255 2.665 ;
        RECT  4.915 2.115 5.250 2.665 ;
        RECT  4.895 3.945 5.125 4.365 ;
        RECT  4.895 0.770 5.120 1.110 ;
        RECT  4.910 2.115 4.915 2.455 ;
        RECT  4.780 0.770 4.895 1.420 ;
        RECT  4.005 3.945 4.895 4.175 ;
        RECT  4.665 0.825 4.780 1.420 ;
        RECT  2.860 1.190 4.665 1.420 ;
        RECT  3.795 2.935 4.005 4.355 ;
        RECT  3.560 1.655 3.900 2.055 ;
        RECT  3.775 2.395 3.795 4.355 ;
        RECT  3.565 2.395 3.775 3.165 ;
        RECT  2.930 4.125 3.775 4.355 ;
        RECT  3.235 2.395 3.565 2.625 ;
        RECT  3.535 1.655 3.560 2.000 ;
        RECT  3.275 3.460 3.460 3.800 ;
        RECT  3.045 2.935 3.275 3.800 ;
        RECT  3.005 1.705 3.235 2.625 ;
        RECT  2.695 2.935 3.045 3.165 ;
        RECT  2.895 1.705 3.005 2.055 ;
        RECT  2.590 4.070 2.930 4.410 ;
        RECT  2.840 1.715 2.895 2.055 ;
        RECT  2.525 0.900 2.860 1.420 ;
        RECT  2.525 2.545 2.695 3.165 ;
        RECT  2.385 4.070 2.590 4.355 ;
        RECT  2.465 0.900 2.525 3.165 ;
        RECT  2.295 0.900 2.465 2.775 ;
        RECT  2.155 3.620 2.385 4.355 ;
        RECT  0.600 3.620 2.155 3.850 ;
        RECT  0.450 3.510 0.600 3.850 ;
        RECT  0.450 1.040 0.560 1.380 ;
        RECT  0.220 1.040 0.450 3.850 ;
    END
END DFFNRXL

MACRO DFFNRX4
    CLASS CORE ;
    FOREIGN DFFNRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNRXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.680 2.745 5.140 3.495 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.960 1.195 18.340 3.220 ;
        RECT  17.940 1.195 17.960 1.535 ;
        RECT  17.940 2.780 17.960 3.120 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.560 1.260 19.660 3.120 ;
        RECT  19.280 1.195 19.560 3.120 ;
        RECT  19.275 1.195 19.280 2.075 ;
        RECT  19.220 2.780 19.280 3.120 ;
        RECT  19.220 1.195 19.275 1.535 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 2.560 1.910 2.900 ;
        RECT  1.460 1.820 1.845 2.900 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.660 2.175 1.180 2.730 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.200 -0.400 20.460 0.400 ;
        RECT  19.860 -0.400 20.200 0.950 ;
        RECT  18.920 -0.400 19.860 0.400 ;
        RECT  18.580 -0.400 18.920 0.950 ;
        RECT  17.640 -0.400 18.580 0.400 ;
        RECT  17.300 -0.400 17.640 0.950 ;
        RECT  16.270 -0.400 17.300 0.400 ;
        RECT  15.930 -0.400 16.270 0.950 ;
        RECT  14.830 -0.400 15.930 0.400 ;
        RECT  14.490 -0.400 14.830 0.950 ;
        RECT  13.370 -0.400 14.490 0.400 ;
        RECT  13.030 -0.400 13.370 0.950 ;
        RECT  11.600 -0.400 13.030 0.400 ;
        RECT  11.260 -0.400 11.600 0.575 ;
        RECT  9.005 -0.400 11.260 0.400 ;
        RECT  8.775 -0.400 9.005 1.475 ;
        RECT  7.150 -0.400 8.775 0.400 ;
        RECT  8.590 1.245 8.775 1.475 ;
        RECT  6.810 -0.400 7.150 0.960 ;
        RECT  5.140 -0.400 6.810 0.400 ;
        RECT  4.800 -0.400 5.140 1.335 ;
        RECT  1.080 -0.400 4.800 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.200 4.640 20.460 5.440 ;
        RECT  19.860 4.040 20.200 5.440 ;
        RECT  18.920 4.640 19.860 5.440 ;
        RECT  18.580 4.040 18.920 5.440 ;
        RECT  17.640 4.640 18.580 5.440 ;
        RECT  17.300 4.040 17.640 5.440 ;
        RECT  16.070 4.640 17.300 5.440 ;
        RECT  15.730 3.055 16.070 5.440 ;
        RECT  13.470 4.640 15.730 5.440 ;
        RECT  13.130 4.080 13.470 5.440 ;
        RECT  10.990 4.640 13.130 5.440 ;
        RECT  10.650 3.675 10.990 5.440 ;
        RECT  8.140 4.640 10.650 5.440 ;
        RECT  7.800 3.920 8.140 5.440 ;
        RECT  4.480 4.640 7.800 5.440 ;
        RECT  4.140 4.465 4.480 5.440 ;
        RECT  1.545 4.640 4.140 5.440 ;
        RECT  1.205 4.465 1.545 5.440 ;
        RECT  0.000 4.640 1.205 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.965 2.030 20.195 3.750 ;
        RECT  17.635 3.520 19.965 3.750 ;
        RECT  17.405 1.395 17.635 3.750 ;
        RECT  16.950 1.395 17.405 1.730 ;
        RECT  16.790 3.265 17.405 3.495 ;
        RECT  16.170 2.100 17.110 2.440 ;
        RECT  16.610 1.390 16.950 1.730 ;
        RECT  16.450 2.975 16.790 3.785 ;
        RECT  16.600 1.395 16.610 1.675 ;
        RECT  15.550 2.155 16.170 2.385 ;
        RECT  15.320 0.720 15.550 2.690 ;
        RECT  15.210 0.720 15.320 1.475 ;
        RECT  14.790 2.460 15.320 2.690 ;
        RECT  14.110 1.245 15.210 1.475 ;
        RECT  14.715 1.725 15.070 2.065 ;
        RECT  14.560 2.460 14.790 3.835 ;
        RECT  14.130 1.725 14.715 2.105 ;
        RECT  14.450 2.985 14.560 3.835 ;
        RECT  12.860 3.605 14.450 3.835 ;
        RECT  13.125 1.875 14.130 2.105 ;
        RECT  13.880 0.700 14.110 1.475 ;
        RECT  13.770 0.700 13.880 1.040 ;
        RECT  12.895 1.495 13.125 3.365 ;
        RECT  10.555 1.495 12.895 1.735 ;
        RECT  12.265 3.135 12.895 3.365 ;
        RECT  12.630 3.605 12.860 4.250 ;
        RECT  12.125 2.425 12.465 2.820 ;
        RECT  11.020 0.955 12.380 1.185 ;
        RECT  12.265 3.750 12.320 4.090 ;
        RECT  12.035 3.135 12.265 4.090 ;
        RECT  10.095 2.425 12.125 2.655 ;
        RECT  10.355 3.135 12.035 3.365 ;
        RECT  11.980 3.750 12.035 4.090 ;
        RECT  10.790 0.635 11.020 1.185 ;
        RECT  9.555 0.635 10.790 0.865 ;
        RECT  10.325 1.095 10.555 1.735 ;
        RECT  10.125 3.135 10.355 3.855 ;
        RECT  9.910 1.095 10.325 1.325 ;
        RECT  9.710 3.625 10.125 3.855 ;
        RECT  9.865 1.720 10.095 2.655 ;
        RECT  9.370 3.625 9.710 3.990 ;
        RECT  9.555 1.745 9.580 3.145 ;
        RECT  9.350 0.635 9.555 3.145 ;
        RECT  9.325 0.635 9.350 1.975 ;
        RECT  9.065 2.915 9.350 3.145 ;
        RECT  8.125 1.715 9.325 1.975 ;
        RECT  7.535 2.205 9.120 2.435 ;
        RECT  8.900 2.915 9.065 3.945 ;
        RECT  8.675 2.915 8.900 4.000 ;
        RECT  8.560 3.660 8.675 4.000 ;
        RECT  8.165 2.840 8.330 3.180 ;
        RECT  7.935 2.840 8.165 3.660 ;
        RECT  7.895 0.675 8.125 1.975 ;
        RECT  7.405 3.430 7.935 3.660 ;
        RECT  7.400 0.675 7.895 0.905 ;
        RECT  7.305 1.565 7.535 3.145 ;
        RECT  7.175 3.430 7.405 4.365 ;
        RECT  6.590 1.565 7.305 1.795 ;
        RECT  6.860 2.915 7.305 3.145 ;
        RECT  5.025 4.135 7.175 4.365 ;
        RECT  6.520 2.915 6.860 3.870 ;
        RECT  6.490 2.100 6.830 2.440 ;
        RECT  6.250 1.430 6.590 1.795 ;
        RECT  5.675 2.155 6.490 2.385 ;
        RECT  4.120 1.565 6.250 1.795 ;
        RECT  5.675 3.560 5.730 3.900 ;
        RECT  5.445 2.025 5.675 3.900 ;
        RECT  4.930 2.025 5.445 2.255 ;
        RECT  5.390 3.560 5.445 3.900 ;
        RECT  4.795 3.945 5.025 4.365 ;
        RECT  3.825 3.945 4.795 4.175 ;
        RECT  4.265 2.320 4.320 2.660 ;
        RECT  2.985 0.825 4.310 1.055 ;
        RECT  4.120 2.245 4.265 2.660 ;
        RECT  3.980 1.565 4.120 2.660 ;
        RECT  3.890 1.565 3.980 2.475 ;
        RECT  3.595 3.035 3.825 4.345 ;
        RECT  3.480 3.035 3.595 3.265 ;
        RECT  2.435 4.115 3.595 4.345 ;
        RECT  3.250 1.980 3.480 3.265 ;
        RECT  3.200 1.980 3.250 2.210 ;
        RECT  2.915 1.820 3.200 2.210 ;
        RECT  3.020 3.500 3.155 3.840 ;
        RECT  2.790 2.465 3.020 3.840 ;
        RECT  2.760 0.825 2.985 1.415 ;
        RECT  2.860 1.820 2.915 2.160 ;
        RECT  2.425 2.465 2.790 2.695 ;
        RECT  2.755 0.825 2.760 1.470 ;
        RECT  2.425 1.130 2.755 1.470 ;
        RECT  2.205 4.005 2.435 4.345 ;
        RECT  2.420 1.130 2.425 2.695 ;
        RECT  2.195 1.185 2.420 2.695 ;
        RECT  0.405 4.005 2.205 4.235 ;
        RECT  0.465 1.220 0.520 1.560 ;
        RECT  0.405 3.180 0.520 3.520 ;
        RECT  0.405 1.215 0.465 1.560 ;
        RECT  0.175 1.215 0.405 4.235 ;
    END
END DFFNRX4

MACRO DFFNRX2
    CLASS CORE ;
    FOREIGN DFFNRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.605 2.875 4.660 3.390 ;
        RECT  4.320 2.755 4.605 3.390 ;
        RECT  4.175 2.755 4.320 3.335 ;
        RECT  4.130 2.875 4.175 3.240 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.565 1.425 15.700 2.100 ;
        RECT  15.565 2.930 15.620 3.270 ;
        RECT  15.335 1.425 15.565 3.270 ;
        RECT  15.280 1.425 15.335 2.100 ;
        RECT  15.280 2.930 15.335 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.705 1.425 17.005 3.270 ;
        RECT  16.590 1.425 16.705 1.765 ;
        RECT  16.570 2.930 16.705 3.270 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 1.550 1.840 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.625 2.480 1.180 3.220 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.265 -0.400 17.160 0.400 ;
        RECT  15.925 -0.400 16.265 1.045 ;
        RECT  14.120 -0.400 15.925 0.400 ;
        RECT  13.780 -0.400 14.120 1.190 ;
        RECT  12.630 -0.400 13.780 0.400 ;
        RECT  12.290 -0.400 12.630 0.575 ;
        RECT  10.540 -0.400 12.290 0.400 ;
        RECT  10.200 -0.400 10.540 0.575 ;
        RECT  8.040 -0.400 10.200 0.400 ;
        RECT  7.700 -0.400 8.040 1.370 ;
        RECT  6.340 -0.400 7.700 0.400 ;
        RECT  6.000 -0.400 6.340 0.960 ;
        RECT  5.120 -0.400 6.000 0.440 ;
        RECT  4.695 -0.400 5.120 1.335 ;
        RECT  1.315 -0.400 4.695 0.400 ;
        RECT  0.975 -0.400 1.315 0.575 ;
        RECT  0.000 -0.400 0.975 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.260 4.640 17.160 5.440 ;
        RECT  15.920 4.080 16.260 5.440 ;
        RECT  14.200 4.640 15.920 5.440 ;
        RECT  13.860 3.680 14.200 5.440 ;
        RECT  11.420 4.640 13.860 5.440 ;
        RECT  11.080 4.080 11.420 5.440 ;
        RECT  8.760 4.640 11.080 5.440 ;
        RECT  7.260 4.080 8.760 5.440 ;
        RECT  4.360 4.640 7.260 5.440 ;
        RECT  4.020 4.465 4.360 5.440 ;
        RECT  1.310 4.640 4.020 5.440 ;
        RECT  0.970 4.465 1.310 5.440 ;
        RECT  0.000 4.640 0.970 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.245 2.095 16.475 2.655 ;
        RECT  16.200 2.425 16.245 2.655 ;
        RECT  15.970 2.425 16.200 3.805 ;
        RECT  14.920 3.575 15.970 3.805 ;
        RECT  14.810 3.575 14.920 4.020 ;
        RECT  14.810 0.850 14.880 1.190 ;
        RECT  14.580 0.850 14.810 4.020 ;
        RECT  14.540 0.850 14.580 1.190 ;
        RECT  14.295 1.590 14.350 2.045 ;
        RECT  14.065 1.590 14.295 3.165 ;
        RECT  14.010 1.590 14.065 2.045 ;
        RECT  13.520 2.935 14.065 3.165 ;
        RECT  13.400 1.815 14.010 2.045 ;
        RECT  13.290 2.935 13.520 3.510 ;
        RECT  13.170 0.910 13.400 2.045 ;
        RECT  12.740 3.280 13.290 3.510 ;
        RECT  13.060 0.910 13.170 1.250 ;
        RECT  12.490 1.815 13.170 2.045 ;
        RECT  12.630 3.280 12.740 3.620 ;
        RECT  12.400 3.280 12.630 4.270 ;
        RECT  12.050 2.460 12.550 2.800 ;
        RECT  12.205 1.630 12.490 2.045 ;
        RECT  12.120 3.930 12.400 4.270 ;
        RECT  12.150 1.630 12.205 1.970 ;
        RECT  11.920 2.460 12.050 3.335 ;
        RECT  11.715 1.685 11.920 3.335 ;
        RECT  11.540 0.635 11.820 0.975 ;
        RECT  11.690 1.270 11.715 3.335 ;
        RECT  11.485 1.270 11.690 1.915 ;
        RECT  11.680 2.680 11.690 3.335 ;
        RECT  10.665 3.105 11.680 3.335 ;
        RECT  11.480 0.635 11.540 1.040 ;
        RECT  9.460 1.270 11.485 1.500 ;
        RECT  11.310 0.690 11.480 1.040 ;
        RECT  11.405 2.205 11.460 2.435 ;
        RECT  11.175 2.205 11.405 2.440 ;
        RECT  9.940 0.810 11.310 1.040 ;
        RECT  10.785 2.210 11.175 2.440 ;
        RECT  10.555 2.040 10.785 2.440 ;
        RECT  10.435 3.105 10.665 3.480 ;
        RECT  9.680 2.040 10.555 2.270 ;
        RECT  10.100 3.250 10.435 3.480 ;
        RECT  9.760 3.250 10.100 3.590 ;
        RECT  9.710 0.630 9.940 1.040 ;
        RECT  9.520 2.600 9.860 2.940 ;
        RECT  8.755 0.630 9.710 0.860 ;
        RECT  9.395 1.735 9.680 2.270 ;
        RECT  9.000 2.655 9.520 2.885 ;
        RECT  9.230 1.090 9.460 1.500 ;
        RECT  9.340 1.735 9.395 2.075 ;
        RECT  9.060 1.090 9.230 1.430 ;
        RECT  8.770 1.705 9.000 3.570 ;
        RECT  8.755 1.705 8.770 1.935 ;
        RECT  7.830 3.205 8.770 3.570 ;
        RECT  8.525 0.630 8.755 1.935 ;
        RECT  8.200 2.170 8.540 2.885 ;
        RECT  7.240 1.705 8.525 1.935 ;
        RECT  6.575 2.170 8.200 2.400 ;
        RECT  7.530 2.630 7.870 2.970 ;
        RECT  7.375 2.740 7.530 2.970 ;
        RECT  7.145 2.740 7.375 3.725 ;
        RECT  7.235 1.205 7.240 1.935 ;
        RECT  7.125 1.150 7.235 1.935 ;
        RECT  6.935 3.495 7.145 3.725 ;
        RECT  6.895 0.665 7.125 1.935 ;
        RECT  6.705 3.495 6.935 4.355 ;
        RECT  6.630 0.665 6.895 0.895 ;
        RECT  4.825 4.125 6.705 4.355 ;
        RECT  6.345 1.575 6.575 3.185 ;
        RECT  5.840 1.575 6.345 1.805 ;
        RECT  6.155 2.955 6.345 3.185 ;
        RECT  6.155 3.470 6.210 3.810 ;
        RECT  5.925 2.955 6.155 3.810 ;
        RECT  5.775 2.140 6.115 2.480 ;
        RECT  5.870 3.470 5.925 3.810 ;
        RECT  5.610 1.455 5.840 1.805 ;
        RECT  5.345 2.195 5.775 2.425 ;
        RECT  5.500 1.455 5.610 1.795 ;
        RECT  3.680 1.565 5.500 1.795 ;
        RECT  5.345 3.550 5.400 3.890 ;
        RECT  5.115 2.195 5.345 3.890 ;
        RECT  5.110 2.195 5.115 2.425 ;
        RECT  5.060 3.550 5.115 3.890 ;
        RECT  4.560 2.030 5.110 2.425 ;
        RECT  4.595 3.945 4.825 4.355 ;
        RECT  3.705 3.945 4.595 4.175 ;
        RECT  4.080 0.675 4.420 1.110 ;
        RECT  2.660 0.675 4.080 0.905 ;
        RECT  3.475 2.395 3.705 4.255 ;
        RECT  3.350 1.565 3.680 2.085 ;
        RECT  2.945 2.395 3.475 2.625 ;
        RECT  2.560 4.025 3.475 4.255 ;
        RECT  3.340 1.745 3.350 2.085 ;
        RECT  2.760 3.300 3.100 3.640 ;
        RECT  2.940 1.655 2.945 2.625 ;
        RECT  2.715 1.600 2.940 2.625 ;
        RECT  2.365 3.300 2.760 3.530 ;
        RECT  2.600 1.600 2.715 1.940 ;
        RECT  2.430 0.675 2.660 1.270 ;
        RECT  2.220 3.970 2.560 4.310 ;
        RECT  2.365 0.905 2.430 1.270 ;
        RECT  2.135 0.905 2.365 3.530 ;
        RECT  0.520 4.005 2.220 4.235 ;
        RECT  0.395 1.060 0.520 1.400 ;
        RECT  0.395 3.520 0.520 4.235 ;
        RECT  0.180 1.060 0.395 4.235 ;
        RECT  0.165 1.100 0.180 4.235 ;
    END
END DFFNRX2

MACRO DFFNRX1
    CLASS CORE ;
    FOREIGN DFFNRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNRXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.525 3.340 4.825 3.570 ;
        RECT  4.130 2.950 4.525 3.570 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.180 2.035 14.410 3.295 ;
        RECT  13.615 2.035 14.180 2.265 ;
        RECT  13.935 3.065 14.180 3.295 ;
        RECT  13.720 3.065 13.935 3.755 ;
        RECT  13.705 3.065 13.720 3.990 ;
        RECT  13.180 3.525 13.705 3.990 ;
        RECT  13.385 1.380 13.615 2.265 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.995 1.355 15.000 1.850 ;
        RECT  14.735 1.260 14.995 3.980 ;
        RECT  14.660 1.260 14.735 1.850 ;
        RECT  14.440 3.640 14.735 3.980 ;
        RECT  14.590 1.260 14.660 1.750 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.730 1.780 2.120 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.680 2.670 1.180 3.220 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.330 -0.400 15.180 0.400 ;
        RECT  13.990 -0.400 14.330 0.575 ;
        RECT  12.250 -0.400 13.990 0.400 ;
        RECT  11.910 -0.400 12.250 0.575 ;
        RECT  10.690 -0.400 11.910 0.400 ;
        RECT  10.350 -0.400 10.690 1.310 ;
        RECT  5.975 -0.400 10.350 0.400 ;
        RECT  7.810 1.440 7.920 1.780 ;
        RECT  7.580 1.205 7.810 1.780 ;
        RECT  6.330 1.205 7.580 1.435 ;
        RECT  5.975 1.205 6.330 1.525 ;
        RECT  5.745 -0.400 5.975 1.525 ;
        RECT  4.020 -0.400 5.745 0.400 ;
        RECT  3.680 -0.400 4.020 0.960 ;
        RECT  1.115 -0.400 3.680 0.400 ;
        RECT  0.775 -0.400 1.115 0.575 ;
        RECT  0.000 -0.400 0.775 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.100 4.640 15.180 5.440 ;
        RECT  13.760 4.465 14.100 5.440 ;
        RECT  12.760 4.640 13.760 5.440 ;
        RECT  12.420 3.620 12.760 5.440 ;
        RECT  10.740 4.640 12.420 5.440 ;
        RECT  10.400 4.070 10.740 5.440 ;
        RECT  8.400 4.640 10.400 5.440 ;
        RECT  7.460 4.070 8.400 5.440 ;
        RECT  4.330 4.640 7.460 5.440 ;
        RECT  3.990 4.465 4.330 5.440 ;
        RECT  1.680 4.640 3.990 5.440 ;
        RECT  1.340 4.465 1.680 5.440 ;
        RECT  0.000 4.640 1.340 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.420 2.495 13.950 2.835 ;
        RECT  13.145 2.495 13.420 3.140 ;
        RECT  13.080 1.250 13.145 3.140 ;
        RECT  12.845 1.250 13.080 2.795 ;
        RECT  12.790 1.250 12.845 1.550 ;
        RECT  12.450 1.210 12.790 1.550 ;
        RECT  12.455 1.825 12.560 2.110 ;
        RECT  12.225 1.825 12.455 3.295 ;
        RECT  11.925 1.825 12.225 2.055 ;
        RECT  11.480 3.065 12.225 3.295 ;
        RECT  11.695 1.595 11.925 2.055 ;
        RECT  11.390 1.595 11.695 1.825 ;
        RECT  11.140 3.065 11.480 3.940 ;
        RECT  11.390 0.970 11.450 1.310 ;
        RECT  11.110 0.970 11.390 1.825 ;
        RECT  11.325 2.140 11.380 2.480 ;
        RECT  11.040 2.140 11.325 2.505 ;
        RECT  10.540 1.595 11.110 1.825 ;
        RECT  9.915 2.275 11.040 2.505 ;
        RECT  10.255 1.595 10.540 2.045 ;
        RECT  10.200 1.705 10.255 2.045 ;
        RECT  9.915 4.000 10.030 4.340 ;
        RECT  9.905 2.275 9.915 4.340 ;
        RECT  9.685 2.020 9.905 4.340 ;
        RECT  9.675 2.020 9.685 4.285 ;
        RECT  9.225 2.020 9.675 2.250 ;
        RECT  9.220 0.650 9.560 0.990 ;
        RECT  9.225 1.230 9.280 1.570 ;
        RECT  8.605 2.500 9.260 2.840 ;
        RECT  8.995 1.230 9.225 2.250 ;
        RECT  8.605 0.675 9.220 0.905 ;
        RECT  8.940 1.230 8.995 1.570 ;
        RECT  8.375 0.675 8.605 3.330 ;
        RECT  6.545 0.675 8.375 0.905 ;
        RECT  8.120 3.100 8.375 3.330 ;
        RECT  7.780 3.100 8.120 3.440 ;
        RECT  8.005 2.020 8.060 2.410 ;
        RECT  7.720 2.020 8.005 2.415 ;
        RECT  6.645 2.180 7.720 2.415 ;
        RECT  7.295 2.705 7.525 3.825 ;
        RECT  7.165 3.595 7.295 3.825 ;
        RECT  6.935 3.595 7.165 4.365 ;
        RECT  4.790 4.135 6.935 4.365 ;
        RECT  6.415 1.825 6.645 3.385 ;
        RECT  6.205 0.635 6.545 0.975 ;
        RECT  5.380 1.825 6.415 2.055 ;
        RECT  6.110 3.155 6.415 3.385 ;
        RECT  5.880 3.155 6.110 3.820 ;
        RECT  5.760 2.440 6.100 2.780 ;
        RECT  5.770 3.480 5.880 3.820 ;
        RECT  5.355 2.495 5.760 2.725 ;
        RECT  5.355 3.480 5.410 3.820 ;
        RECT  5.370 1.655 5.380 2.055 ;
        RECT  5.150 1.180 5.370 2.055 ;
        RECT  5.125 2.435 5.355 3.820 ;
        RECT  5.140 1.180 5.150 1.885 ;
        RECT  3.570 1.655 5.140 1.885 ;
        RECT  4.920 2.435 5.125 2.665 ;
        RECT  5.070 3.480 5.125 3.820 ;
        RECT  4.555 2.120 4.920 2.665 ;
        RECT  4.565 0.770 4.870 1.110 ;
        RECT  4.560 3.945 4.790 4.365 ;
        RECT  4.335 0.770 4.565 1.420 ;
        RECT  3.675 3.945 4.560 4.175 ;
        RECT  2.530 1.190 4.335 1.420 ;
        RECT  3.465 2.935 3.675 4.355 ;
        RECT  3.230 1.655 3.570 2.080 ;
        RECT  3.445 2.395 3.465 4.355 ;
        RECT  3.235 2.395 3.445 3.165 ;
        RECT  2.145 4.125 3.445 4.355 ;
        RECT  2.905 2.395 3.235 2.625 ;
        RECT  2.775 3.480 3.110 3.840 ;
        RECT  2.845 2.105 2.905 2.625 ;
        RECT  2.675 1.940 2.845 2.625 ;
        RECT  2.545 2.855 2.775 3.840 ;
        RECT  2.615 1.940 2.675 2.335 ;
        RECT  2.380 2.855 2.545 3.085 ;
        RECT  2.380 1.160 2.530 1.500 ;
        RECT  2.190 1.160 2.380 3.085 ;
        RECT  2.150 1.220 2.190 3.085 ;
        RECT  1.915 3.745 2.145 4.355 ;
        RECT  0.845 3.745 1.915 3.975 ;
        RECT  0.505 3.520 0.845 3.975 ;
        RECT  0.390 1.150 0.520 1.490 ;
        RECT  0.390 3.520 0.505 3.750 ;
        RECT  0.180 1.150 0.390 3.750 ;
        RECT  0.160 1.260 0.180 3.750 ;
    END
END DFFNRX1

MACRO DFFNXL
    CLASS CORE ;
    FOREIGN DFFNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 1.200 11.040 3.790 ;
        RECT  10.600 3.450 10.700 3.790 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 0.865 10.345 3.420 ;
        RECT  10.040 0.865 10.115 1.285 ;
        RECT  9.290 3.190 10.115 3.420 ;
        RECT  9.830 0.865 10.040 1.095 ;
        RECT  9.300 0.745 9.830 1.095 ;
        RECT  8.950 3.190 9.290 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 1.675 1.840 2.320 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.630 1.180 3.220 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.460 -0.400 11.220 0.400 ;
        RECT  10.120 -0.400 10.460 0.575 ;
        RECT  8.880 -0.400 10.120 0.400 ;
        RECT  8.540 -0.400 8.880 0.575 ;
        RECT  6.400 -0.400 8.540 0.400 ;
        RECT  6.060 -0.400 6.400 1.555 ;
        RECT  4.070 -0.400 6.060 0.400 ;
        RECT  3.730 -0.400 4.070 1.150 ;
        RECT  1.265 -0.400 3.730 0.400 ;
        RECT  0.925 -0.400 1.265 0.575 ;
        RECT  0.000 -0.400 0.925 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.180 4.640 11.220 5.440 ;
        RECT  9.840 4.410 10.180 5.440 ;
        RECT  8.470 4.640 9.840 5.440 ;
        RECT  8.130 4.465 8.470 5.440 ;
        RECT  5.795 4.640 8.130 5.440 ;
        RECT  5.455 4.465 5.795 5.440 ;
        RECT  1.485 4.640 5.455 5.440 ;
        RECT  1.145 4.410 1.485 5.440 ;
        RECT  0.000 4.640 1.145 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.805 2.005 9.870 2.375 ;
        RECT  9.680 1.470 9.805 2.945 ;
        RECT  9.575 1.460 9.680 2.945 ;
        RECT  9.340 1.460 9.575 1.800 ;
        RECT  8.400 2.715 9.575 2.945 ;
        RECT  8.915 2.105 9.255 2.445 ;
        RECT  9.175 4.060 9.230 4.400 ;
        RECT  8.890 3.970 9.175 4.400 ;
        RECT  8.880 2.105 8.915 2.335 ;
        RECT  8.400 3.970 8.890 4.200 ;
        RECT  8.650 1.440 8.880 2.335 ;
        RECT  7.550 1.440 8.650 1.835 ;
        RECT  8.350 2.715 8.400 4.200 ;
        RECT  8.170 2.180 8.350 4.200 ;
        RECT  8.010 2.180 8.170 2.945 ;
        RECT  7.760 0.835 8.100 1.175 ;
        RECT  6.940 0.945 7.760 1.175 ;
        RECT  7.320 1.440 7.550 4.150 ;
        RECT  7.260 3.920 7.320 4.150 ;
        RECT  6.920 3.920 7.260 4.260 ;
        RECT  6.980 1.840 7.090 3.160 ;
        RECT  6.940 1.840 6.980 3.615 ;
        RECT  6.750 0.945 6.940 3.615 ;
        RECT  6.710 0.945 6.750 2.070 ;
        RECT  6.270 3.385 6.750 3.615 ;
        RECT  5.600 1.840 6.710 2.070 ;
        RECT  6.310 2.380 6.420 2.720 ;
        RECT  6.080 2.380 6.310 3.135 ;
        RECT  6.040 3.385 6.270 4.235 ;
        RECT  5.800 2.905 6.080 3.135 ;
        RECT  3.590 4.005 6.040 4.235 ;
        RECT  5.570 2.905 5.800 3.775 ;
        RECT  5.330 1.210 5.600 2.070 ;
        RECT  4.760 3.545 5.570 3.775 ;
        RECT  5.260 1.210 5.330 3.120 ;
        RECT  5.100 1.840 5.260 3.120 ;
        RECT  4.990 2.780 5.100 3.120 ;
        RECT  4.815 0.830 4.870 1.170 ;
        RECT  4.760 0.830 4.815 2.470 ;
        RECT  4.585 0.830 4.760 3.775 ;
        RECT  4.530 0.830 4.585 1.170 ;
        RECT  4.490 2.220 4.585 3.775 ;
        RECT  3.580 2.220 4.490 2.560 ;
        RECT  4.015 1.485 4.355 1.825 ;
        RECT  3.375 1.595 4.015 1.825 ;
        RECT  3.480 3.950 3.590 4.290 ;
        RECT  3.250 3.720 3.480 4.290 ;
        RECT  3.295 1.195 3.375 1.825 ;
        RECT  3.295 3.150 3.350 3.490 ;
        RECT  3.065 1.195 3.295 3.490 ;
        RECT  2.490 3.720 3.250 3.950 ;
        RECT  2.710 1.195 3.065 1.480 ;
        RECT  3.010 3.150 3.065 3.490 ;
        RECT  2.030 4.180 2.895 4.410 ;
        RECT  2.370 1.140 2.710 1.480 ;
        RECT  2.430 1.845 2.490 3.950 ;
        RECT  2.260 1.735 2.430 3.950 ;
        RECT  2.090 1.735 2.260 2.075 ;
        RECT  1.800 3.605 2.030 4.410 ;
        RECT  0.650 3.605 1.800 3.835 ;
        RECT  0.415 3.455 0.650 3.835 ;
        RECT  0.415 1.200 0.530 1.540 ;
        RECT  0.190 1.200 0.415 3.835 ;
        RECT  0.185 1.255 0.190 3.835 ;
    END
END DFFNXL

MACRO DFFNX4
    CLASS CORE ;
    FOREIGN DFFNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.010 1.820 15.040 3.220 ;
        RECT  14.965 1.290 15.010 3.220 ;
        RECT  14.945 1.290 14.965 3.225 ;
        RECT  14.670 1.290 14.945 3.280 ;
        RECT  14.660 1.820 14.670 3.280 ;
        RECT  14.605 2.940 14.660 3.280 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.720 1.290 13.730 1.850 ;
        RECT  13.675 1.290 13.720 3.220 ;
        RECT  13.665 1.290 13.675 3.225 ;
        RECT  13.390 1.290 13.665 3.280 ;
        RECT  13.340 1.820 13.390 3.280 ;
        RECT  13.325 2.940 13.340 3.280 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.365 2.400 1.595 3.185 ;
        RECT  1.125 2.890 1.365 3.185 ;
        RECT  1.105 2.955 1.125 3.185 ;
        RECT  0.875 2.955 1.105 3.195 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 1.845 1.765 2.075 ;
        RECT  0.695 1.845 0.925 2.250 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.650 -0.400 15.840 0.400 ;
        RECT  15.310 -0.400 15.650 0.965 ;
        RECT  14.370 -0.400 15.310 0.400 ;
        RECT  14.030 -0.400 14.370 0.965 ;
        RECT  13.090 -0.400 14.030 0.400 ;
        RECT  12.750 -0.400 13.090 0.965 ;
        RECT  11.610 -0.400 12.750 0.400 ;
        RECT  11.270 -0.400 11.610 0.575 ;
        RECT  8.910 -0.400 11.270 0.400 ;
        RECT  8.570 -0.400 8.910 1.280 ;
        RECT  6.350 -0.400 8.570 0.400 ;
        RECT  6.010 -0.400 6.350 1.435 ;
        RECT  3.925 -0.400 6.010 0.400 ;
        RECT  3.585 -0.400 3.925 1.375 ;
        RECT  1.320 -0.400 3.585 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.585 4.640 15.840 5.440 ;
        RECT  15.245 4.075 15.585 5.440 ;
        RECT  14.305 4.640 15.245 5.440 ;
        RECT  13.965 4.075 14.305 5.440 ;
        RECT  13.025 4.640 13.965 5.440 ;
        RECT  12.685 4.075 13.025 5.440 ;
        RECT  11.460 4.640 12.685 5.440 ;
        RECT  11.090 4.400 11.460 5.440 ;
        RECT  8.880 4.640 11.090 5.440 ;
        RECT  8.540 4.090 8.880 5.440 ;
        RECT  6.265 4.640 8.540 5.440 ;
        RECT  5.925 4.465 6.265 5.440 ;
        RECT  4.000 4.640 5.925 5.440 ;
        RECT  3.660 4.465 4.000 5.440 ;
        RECT  1.400 4.640 3.660 5.440 ;
        RECT  1.060 4.465 1.400 5.440 ;
        RECT  0.000 4.640 1.060 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.325 2.290 15.555 3.755 ;
        RECT  12.995 3.525 15.325 3.755 ;
        RECT  12.765 1.265 12.995 3.755 ;
        RECT  12.370 1.265 12.765 1.495 ;
        RECT  12.240 3.420 12.765 3.755 ;
        RECT  12.285 2.290 12.515 3.045 ;
        RECT  12.030 1.130 12.370 1.495 ;
        RECT  10.970 2.815 12.285 3.045 ;
        RECT  11.900 3.420 12.240 3.760 ;
        RECT  11.430 1.265 12.030 1.495 ;
        RECT  11.200 1.265 11.430 2.580 ;
        RECT  10.740 0.995 10.970 3.855 ;
        RECT  9.625 0.995 10.740 1.225 ;
        RECT  10.160 3.625 10.740 3.855 ;
        RECT  10.275 1.495 10.505 2.905 ;
        RECT  9.920 2.675 10.275 2.905 ;
        RECT  9.820 3.625 10.160 3.990 ;
        RECT  9.810 2.595 9.920 2.935 ;
        RECT  7.600 3.625 9.820 3.855 ;
        RECT  9.580 2.595 9.810 3.335 ;
        RECT  9.395 0.995 9.625 1.825 ;
        RECT  7.590 3.105 9.580 3.335 ;
        RECT  7.685 1.595 9.395 1.825 ;
        RECT  8.820 2.140 9.110 2.480 ;
        RECT  8.300 2.065 8.820 2.480 ;
        RECT  6.615 2.065 8.300 2.295 ;
        RECT  7.630 1.330 7.685 1.825 ;
        RECT  7.455 1.275 7.630 1.825 ;
        RECT  7.315 3.625 7.600 4.080 ;
        RECT  7.250 2.530 7.590 3.335 ;
        RECT  7.290 1.275 7.455 1.615 ;
        RECT  7.260 3.740 7.315 4.080 ;
        RECT  5.480 3.105 7.250 3.335 ;
        RECT  6.205 1.670 6.615 2.360 ;
        RECT  5.780 1.670 6.205 1.900 ;
        RECT  5.550 0.935 5.780 1.900 ;
        RECT  4.685 0.935 5.550 1.165 ;
        RECT  5.425 3.060 5.480 3.400 ;
        RECT  5.320 3.060 5.425 4.175 ;
        RECT  5.195 1.420 5.320 4.175 ;
        RECT  5.090 1.420 5.195 3.425 ;
        RECT  3.205 3.945 5.195 4.175 ;
        RECT  4.685 2.720 4.705 3.710 ;
        RECT  4.475 0.935 4.685 3.710 ;
        RECT  4.455 0.935 4.475 2.950 ;
        RECT  4.310 1.130 4.455 1.470 ;
        RECT  3.365 2.610 4.455 2.950 ;
        RECT  3.800 1.890 4.140 2.230 ;
        RECT  3.095 1.945 3.800 2.175 ;
        RECT  2.975 3.945 3.205 4.235 ;
        RECT  3.065 1.375 3.095 2.175 ;
        RECT  2.835 1.375 3.065 3.515 ;
        RECT  2.165 4.005 2.975 4.235 ;
        RECT  1.780 0.675 2.970 0.905 ;
        RECT  2.540 1.375 2.835 1.605 ;
        RECT  2.665 3.285 2.835 3.515 ;
        RECT  2.435 3.285 2.665 3.650 ;
        RECT  2.255 1.240 2.540 1.605 ;
        RECT  2.165 1.920 2.305 2.995 ;
        RECT  2.200 1.240 2.255 1.580 ;
        RECT  2.075 1.920 2.165 4.235 ;
        RECT  1.935 2.765 2.075 4.235 ;
        RECT  1.550 0.675 1.780 1.395 ;
        RECT  0.560 1.165 1.550 1.395 ;
        RECT  0.430 1.165 0.560 1.530 ;
        RECT  0.430 2.900 0.540 4.180 ;
        RECT  0.275 1.165 0.430 4.180 ;
        RECT  0.220 1.190 0.275 4.180 ;
        RECT  0.200 1.245 0.220 4.180 ;
    END
END DFFNX4

MACRO DFFNX2
    CLASS CORE ;
    FOREIGN DFFNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 1.355 12.985 3.330 ;
        RECT  12.680 1.355 12.755 1.845 ;
        RECT  12.700 3.100 12.755 3.330 ;
        RECT  12.360 3.100 12.700 3.440 ;
        RECT  12.580 1.355 12.680 1.695 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.505 0.700 11.560 1.040 ;
        RECT  11.220 0.700 11.505 1.080 ;
        RECT  10.865 0.850 11.220 1.080 ;
        RECT  11.080 2.880 11.160 3.220 ;
        RECT  10.865 2.635 11.080 3.220 ;
        RECT  10.700 0.850 10.865 3.220 ;
        RECT  10.635 0.850 10.700 3.165 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.405 1.825 2.240 ;
        RECT  1.325 1.405 1.460 1.745 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.060 1.180 2.660 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.480 -0.400 13.860 0.400 ;
        RECT  13.140 -0.400 13.480 0.575 ;
        RECT  12.360 -0.400 13.140 0.400 ;
        RECT  12.020 -0.400 12.360 0.575 ;
        RECT  10.760 -0.400 12.020 0.400 ;
        RECT  10.420 -0.400 10.760 0.575 ;
        RECT  8.800 -0.400 10.420 0.400 ;
        RECT  8.460 -0.400 8.800 1.270 ;
        RECT  6.185 -0.400 8.460 0.400 ;
        RECT  5.845 -0.400 6.185 1.440 ;
        RECT  4.020 -0.400 5.845 0.400 ;
        RECT  3.680 -0.400 4.020 1.285 ;
        RECT  1.285 -0.400 3.680 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.260 4.640 13.860 5.440 ;
        RECT  12.920 4.465 13.260 5.440 ;
        RECT  11.920 4.640 12.920 5.440 ;
        RECT  11.580 4.465 11.920 5.440 ;
        RECT  9.940 4.640 11.580 5.440 ;
        RECT  8.190 4.465 9.940 5.440 ;
        RECT  5.870 4.640 8.190 5.440 ;
        RECT  5.530 4.465 5.870 5.440 ;
        RECT  4.530 4.640 5.530 5.440 ;
        RECT  4.190 4.465 4.530 5.440 ;
        RECT  1.340 4.640 4.190 5.440 ;
        RECT  1.000 4.410 1.340 5.440 ;
        RECT  0.000 4.640 1.000 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.435 4.020 12.490 4.360 ;
        RECT  12.150 3.995 12.435 4.360 ;
        RECT  12.125 3.995 12.150 4.225 ;
        RECT  11.895 1.535 12.125 4.225 ;
        RECT  11.220 1.535 11.895 1.765 ;
        RECT  11.160 3.995 11.895 4.225 ;
        RECT  11.435 2.275 11.665 3.680 ;
        RECT  9.975 3.450 11.435 3.680 ;
        RECT  11.050 3.995 11.160 4.370 ;
        RECT  10.820 3.910 11.050 4.370 ;
        RECT  9.640 3.910 10.820 4.140 ;
        RECT  9.745 1.775 9.975 3.680 ;
        RECT  9.600 1.775 9.745 2.005 ;
        RECT  9.030 3.415 9.745 3.680 ;
        RECT  9.370 1.145 9.600 2.005 ;
        RECT  9.110 2.350 9.450 2.690 ;
        RECT  9.260 1.145 9.370 1.795 ;
        RECT  8.130 1.565 9.260 1.795 ;
        RECT  8.195 2.405 9.110 2.635 ;
        RECT  8.920 3.360 9.030 3.700 ;
        RECT  8.690 3.360 8.920 3.960 ;
        RECT  7.155 3.730 8.690 3.960 ;
        RECT  7.965 2.405 8.195 3.130 ;
        RECT  7.900 1.160 8.130 1.795 ;
        RECT  7.300 2.900 7.965 3.130 ;
        RECT  7.520 1.160 7.900 1.390 ;
        RECT  7.180 1.050 7.520 1.390 ;
        RECT  7.210 2.820 7.300 3.160 ;
        RECT  6.980 1.770 7.210 3.160 ;
        RECT  6.925 3.440 7.155 4.275 ;
        RECT  5.390 1.770 6.980 2.000 ;
        RECT  6.960 2.820 6.980 3.160 ;
        RECT  6.330 2.930 6.960 3.160 ;
        RECT  5.860 2.245 6.610 2.475 ;
        RECT  6.100 2.930 6.330 4.235 ;
        RECT  3.595 4.005 6.100 4.235 ;
        RECT  5.630 2.245 5.860 3.755 ;
        RECT  4.695 3.525 5.630 3.755 ;
        RECT  5.390 1.095 5.445 1.435 ;
        RECT  5.380 1.095 5.390 2.000 ;
        RECT  5.330 1.095 5.380 2.910 ;
        RECT  5.150 1.095 5.330 2.965 ;
        RECT  5.105 1.095 5.150 1.435 ;
        RECT  4.990 2.625 5.150 2.965 ;
        RECT  4.685 2.270 4.695 3.755 ;
        RECT  4.465 0.965 4.685 3.755 ;
        RECT  4.455 0.965 4.465 2.580 ;
        RECT  3.925 2.170 4.455 2.500 ;
        RECT  3.355 1.555 4.180 1.785 ;
        RECT  3.585 2.170 3.925 2.510 ;
        RECT  3.365 3.695 3.595 4.235 ;
        RECT  2.895 3.695 3.365 3.925 ;
        RECT  3.125 1.545 3.355 3.430 ;
        RECT  2.970 1.545 3.125 1.785 ;
        RECT  2.740 0.920 2.970 1.785 ;
        RECT  2.665 2.820 2.895 3.925 ;
        RECT  1.980 4.180 2.840 4.410 ;
        RECT  2.660 0.920 2.740 1.150 ;
        RECT  2.375 2.820 2.665 3.050 ;
        RECT  2.320 0.810 2.660 1.150 ;
        RECT  2.375 1.380 2.430 1.720 ;
        RECT  2.145 1.380 2.375 3.050 ;
        RECT  2.090 1.380 2.145 1.720 ;
        RECT  1.750 3.605 1.980 4.410 ;
        RECT  0.790 3.605 1.750 3.835 ;
        RECT  0.570 3.020 0.790 3.835 ;
        RECT  0.390 1.340 0.570 3.835 ;
        RECT  0.340 1.340 0.390 3.310 ;
        RECT  0.180 1.340 0.340 1.680 ;
    END
END DFFNX2

MACRO DFFNX1
    CLASS CORE ;
    FOREIGN DFFNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 1.190 11.040 3.880 ;
        RECT  10.600 3.540 10.700 3.880 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 0.865 10.345 3.420 ;
        RECT  9.640 0.865 10.115 1.095 ;
        RECT  9.230 3.190 10.115 3.420 ;
        RECT  9.300 0.690 9.640 1.095 ;
        RECT  8.890 3.190 9.230 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.820 1.840 2.410 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.685 1.180 3.220 ;
        END
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.460 -0.400 11.220 0.400 ;
        RECT  10.120 -0.400 10.460 0.575 ;
        RECT  8.880 -0.400 10.120 0.400 ;
        RECT  8.540 -0.400 8.880 0.575 ;
        RECT  6.440 -0.400 8.540 0.400 ;
        RECT  6.100 -0.400 6.440 1.460 ;
        RECT  4.070 -0.400 6.100 0.400 ;
        RECT  3.730 -0.400 4.070 1.150 ;
        RECT  1.305 -0.400 3.730 0.400 ;
        RECT  0.965 -0.400 1.305 0.575 ;
        RECT  0.000 -0.400 0.965 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.180 4.640 11.220 5.440 ;
        RECT  9.840 4.410 10.180 5.440 ;
        RECT  8.470 4.640 9.840 5.440 ;
        RECT  8.130 4.465 8.470 5.440 ;
        RECT  5.800 4.640 8.130 5.440 ;
        RECT  4.520 4.465 5.800 5.440 ;
        RECT  1.035 4.640 4.520 5.440 ;
        RECT  0.695 4.410 1.035 5.440 ;
        RECT  0.000 4.640 0.695 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.640 1.470 9.870 2.760 ;
        RECT  9.340 1.470 9.640 1.810 ;
        RECT  8.400 2.530 9.640 2.760 ;
        RECT  8.880 2.065 9.255 2.295 ;
        RECT  8.890 3.990 9.230 4.370 ;
        RECT  8.400 3.990 8.890 4.220 ;
        RECT  8.650 1.440 8.880 2.295 ;
        RECT  7.550 1.440 8.650 1.835 ;
        RECT  8.350 2.530 8.400 4.220 ;
        RECT  8.170 2.180 8.350 4.220 ;
        RECT  8.065 2.180 8.170 2.760 ;
        RECT  6.940 0.670 8.100 0.900 ;
        RECT  8.010 2.180 8.065 2.520 ;
        RECT  7.320 1.440 7.550 4.230 ;
        RECT  7.210 4.000 7.320 4.230 ;
        RECT  6.870 4.000 7.210 4.340 ;
        RECT  6.865 2.820 7.090 3.160 ;
        RECT  6.865 0.670 6.940 1.995 ;
        RECT  6.710 0.670 6.865 3.615 ;
        RECT  6.635 1.765 6.710 3.615 ;
        RECT  5.555 1.840 6.635 2.070 ;
        RECT  6.270 3.385 6.635 3.615 ;
        RECT  6.135 2.380 6.365 3.135 ;
        RECT  6.040 3.385 6.270 4.235 ;
        RECT  5.800 2.905 6.135 3.135 ;
        RECT  3.590 4.005 6.040 4.235 ;
        RECT  5.570 2.905 5.800 3.775 ;
        RECT  5.555 1.170 5.610 1.510 ;
        RECT  4.760 3.545 5.570 3.775 ;
        RECT  5.315 1.170 5.555 2.070 ;
        RECT  5.315 2.790 5.330 3.130 ;
        RECT  5.270 1.170 5.315 3.130 ;
        RECT  5.085 1.840 5.270 3.130 ;
        RECT  4.990 2.790 5.085 3.130 ;
        RECT  4.815 0.830 4.870 1.170 ;
        RECT  4.760 0.830 4.815 2.470 ;
        RECT  4.585 0.830 4.760 3.775 ;
        RECT  4.530 0.830 4.585 1.170 ;
        RECT  4.490 2.200 4.585 3.775 ;
        RECT  3.580 2.200 4.490 2.540 ;
        RECT  4.015 1.425 4.355 1.765 ;
        RECT  3.295 1.425 4.015 1.655 ;
        RECT  3.485 3.950 3.590 4.290 ;
        RECT  3.250 3.720 3.485 4.290 ;
        RECT  3.295 3.150 3.350 3.490 ;
        RECT  3.065 1.170 3.295 3.490 ;
        RECT  2.375 3.720 3.250 3.950 ;
        RECT  2.710 1.170 3.065 1.400 ;
        RECT  3.010 3.150 3.065 3.490 ;
        RECT  1.765 4.180 2.895 4.410 ;
        RECT  2.370 1.060 2.710 1.400 ;
        RECT  2.145 1.685 2.375 3.950 ;
        RECT  1.535 3.605 1.765 4.410 ;
        RECT  0.650 3.605 1.535 3.835 ;
        RECT  0.415 3.455 0.650 3.835 ;
        RECT  0.415 1.095 0.530 1.435 ;
        RECT  0.190 1.095 0.415 3.835 ;
        RECT  0.185 1.150 0.190 3.835 ;
    END
END DFFNX1

MACRO DFFHQXL
    CLASS CORE ;
    FOREIGN DFFHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 0.740 10.435 3.530 ;
        RECT  10.205 0.740 10.345 3.755 ;
        RECT  9.590 0.740 10.205 0.970 ;
        RECT  10.115 3.190 10.205 3.755 ;
        RECT  9.050 3.190 10.115 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 1.820 1.840 2.630 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 2.080 1.105 2.770 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 -0.400 10.560 0.400 ;
        RECT  8.830 -0.400 9.170 0.575 ;
        RECT  6.315 -0.400 8.830 0.400 ;
        RECT  6.085 -0.400 6.315 1.460 ;
        RECT  4.015 -0.400 6.085 0.400 ;
        RECT  3.785 -0.400 4.015 1.150 ;
        RECT  1.350 -0.400 3.785 0.400 ;
        RECT  1.010 -0.400 1.350 0.575 ;
        RECT  0.000 -0.400 1.010 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.630 4.640 10.560 5.440 ;
        RECT  8.290 4.465 8.630 5.440 ;
        RECT  5.795 4.640 8.290 5.440 ;
        RECT  5.455 4.465 5.795 5.440 ;
        RECT  1.815 4.640 5.455 5.440 ;
        RECT  1.475 4.465 1.815 5.440 ;
        RECT  0.000 4.640 1.475 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.925 1.460 9.970 1.800 ;
        RECT  9.695 1.460 9.925 2.960 ;
        RECT  9.630 1.460 9.695 1.800 ;
        RECT  8.640 2.730 9.695 2.960 ;
        RECT  9.235 2.040 9.465 2.380 ;
        RECT  9.090 4.115 9.390 4.345 ;
        RECT  9.170 2.040 9.235 2.270 ;
        RECT  8.940 1.605 9.170 2.270 ;
        RECT  8.860 4.005 9.090 4.345 ;
        RECT  7.955 1.605 8.940 1.835 ;
        RECT  8.640 4.005 8.860 4.235 ;
        RECT  8.410 2.180 8.640 4.235 ;
        RECT  8.300 2.180 8.410 2.520 ;
        RECT  6.775 0.875 8.390 1.105 ;
        RECT  7.725 1.370 7.955 4.375 ;
        RECT  7.030 4.145 7.725 4.375 ;
        RECT  7.265 1.715 7.495 3.915 ;
        RECT  7.235 1.715 7.265 1.945 ;
        RECT  6.595 3.685 7.265 3.915 ;
        RECT  7.005 1.345 7.235 1.945 ;
        RECT  6.805 2.225 7.035 3.455 ;
        RECT  6.775 2.225 6.805 2.455 ;
        RECT  6.135 3.225 6.805 3.455 ;
        RECT  6.545 0.875 6.775 2.455 ;
        RECT  6.365 3.685 6.595 4.140 ;
        RECT  5.560 1.765 6.545 1.995 ;
        RECT  5.675 2.745 6.420 2.975 ;
        RECT  5.905 3.225 6.135 4.235 ;
        RECT  2.375 4.005 5.905 4.235 ;
        RECT  5.445 2.745 5.675 3.775 ;
        RECT  5.365 1.170 5.570 1.510 ;
        RECT  4.680 3.545 5.445 3.775 ;
        RECT  5.275 0.630 5.365 1.510 ;
        RECT  5.215 0.630 5.275 1.940 ;
        RECT  5.135 0.630 5.215 3.130 ;
        RECT  5.045 1.225 5.135 3.130 ;
        RECT  4.985 1.710 5.045 3.130 ;
        RECT  4.680 0.810 4.815 1.465 ;
        RECT  4.585 0.810 4.680 3.775 ;
        RECT  4.450 1.235 4.585 3.775 ;
        RECT  4.395 2.185 4.450 3.775 ;
        RECT  3.920 2.185 4.395 2.415 ;
        RECT  3.295 1.515 4.220 1.745 ;
        RECT  3.580 2.130 3.920 2.470 ;
        RECT  3.065 0.805 3.295 3.680 ;
        RECT  2.370 0.805 3.065 1.035 ;
        RECT  2.145 1.410 2.375 4.235 ;
        RECT  1.055 3.135 2.145 3.365 ;
        RECT  0.715 3.025 1.055 3.365 ;
        RECT  0.415 1.410 0.750 1.750 ;
        RECT  0.415 3.025 0.715 3.255 ;
        RECT  0.185 1.410 0.415 3.255 ;
    END
END DFFHQXL

MACRO DFFHQX4
    CLASS CORE ;
    FOREIGN DFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFHQXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.620 1.820 13.720 3.220 ;
        RECT  13.540 0.835 13.620 3.220 ;
        RECT  13.340 0.835 13.540 3.675 ;
        RECT  13.280 0.835 13.340 1.645 ;
        RECT  13.200 2.865 13.340 3.675 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.415 2.605 1.840 3.280 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 2.200 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.340 -0.400 14.520 0.400 ;
        RECT  14.000 -0.400 14.340 1.015 ;
        RECT  12.860 -0.400 14.000 0.400 ;
        RECT  12.520 -0.400 12.860 0.575 ;
        RECT  11.560 -0.400 12.520 0.400 ;
        RECT  11.220 -0.400 11.560 1.250 ;
        RECT  9.345 -0.400 11.220 0.400 ;
        RECT  9.115 -0.400 9.345 1.270 ;
        RECT  6.205 -0.400 9.115 0.400 ;
        RECT  5.975 -0.400 6.205 1.370 ;
        RECT  3.820 -0.400 5.975 0.400 ;
        RECT  3.480 -0.400 3.820 1.270 ;
        RECT  1.300 -0.400 3.480 0.400 ;
        RECT  0.960 -0.400 1.300 0.575 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.300 4.640 14.520 5.440 ;
        RECT  13.960 4.465 14.300 5.440 ;
        RECT  12.780 4.640 13.960 5.440 ;
        RECT  12.440 4.465 12.780 5.440 ;
        RECT  11.400 4.640 12.440 5.440 ;
        RECT  9.650 4.465 11.400 5.440 ;
        RECT  6.130 4.640 9.650 5.440 ;
        RECT  5.790 4.465 6.130 5.440 ;
        RECT  4.065 4.640 5.790 5.440 ;
        RECT  3.725 4.465 4.065 5.440 ;
        RECT  1.370 4.640 3.725 5.440 ;
        RECT  1.030 4.465 1.370 5.440 ;
        RECT  0.000 4.640 1.030 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.305 2.065 12.310 3.810 ;
        RECT  12.080 1.195 12.305 3.810 ;
        RECT  12.075 1.195 12.080 2.430 ;
        RECT  11.820 3.470 12.080 3.810 ;
        RECT  11.385 2.200 12.075 2.430 ;
        RECT  11.155 2.870 11.840 3.100 ;
        RECT  10.925 1.500 11.155 3.965 ;
        RECT  10.200 1.500 10.925 1.730 ;
        RECT  10.125 3.735 10.925 3.965 ;
        RECT  10.465 1.960 10.695 3.235 ;
        RECT  8.420 1.960 10.465 2.190 ;
        RECT  9.660 3.005 10.465 3.235 ;
        RECT  10.005 2.425 10.235 2.770 ;
        RECT  9.860 0.965 10.200 1.730 ;
        RECT  9.895 3.735 10.125 4.030 ;
        RECT  9.200 2.540 10.005 2.770 ;
        RECT  7.830 3.800 9.895 4.030 ;
        RECT  9.855 1.075 9.860 1.730 ;
        RECT  8.885 1.500 9.855 1.730 ;
        RECT  9.430 3.005 9.660 3.570 ;
        RECT  6.770 3.340 9.430 3.570 ;
        RECT  8.970 2.540 9.200 3.110 ;
        RECT  7.500 2.880 8.970 3.110 ;
        RECT  8.655 1.050 8.885 1.730 ;
        RECT  7.960 2.420 8.740 2.650 ;
        RECT  7.360 1.050 8.655 1.280 ;
        RECT  8.190 1.515 8.420 2.190 ;
        RECT  7.125 1.515 8.190 1.745 ;
        RECT  7.730 2.035 7.960 2.650 ;
        RECT  7.490 3.800 7.830 4.140 ;
        RECT  6.630 2.035 7.730 2.265 ;
        RECT  7.215 2.540 7.500 3.110 ;
        RECT  7.160 2.540 7.215 3.000 ;
        RECT  6.515 2.760 7.160 3.000 ;
        RECT  6.895 1.085 7.125 1.745 ;
        RECT  6.640 1.085 6.895 1.315 ;
        RECT  6.575 2.035 6.630 2.400 ;
        RECT  6.345 1.600 6.575 2.400 ;
        RECT  6.285 2.760 6.515 4.225 ;
        RECT  5.745 1.600 6.345 1.830 ;
        RECT  6.290 2.060 6.345 2.400 ;
        RECT  6.055 2.760 6.285 2.990 ;
        RECT  2.430 3.995 6.285 4.225 ;
        RECT  5.960 2.225 6.055 2.990 ;
        RECT  5.825 2.115 5.960 2.990 ;
        RECT  5.620 2.115 5.825 2.455 ;
        RECT  5.515 0.630 5.745 1.830 ;
        RECT  5.590 3.315 5.720 3.655 ;
        RECT  5.380 2.705 5.590 3.655 ;
        RECT  4.430 0.630 5.515 0.860 ;
        RECT  5.360 2.705 5.380 3.600 ;
        RECT  5.085 2.705 5.360 2.935 ;
        RECT  5.085 1.130 5.285 1.690 ;
        RECT  5.055 1.130 5.085 2.935 ;
        RECT  4.855 1.460 5.055 2.935 ;
        RECT  4.525 3.320 4.865 3.660 ;
        RECT  4.745 1.905 4.855 2.245 ;
        RECT  4.515 1.145 4.540 1.485 ;
        RECT  4.520 3.320 4.525 3.605 ;
        RECT  4.515 2.625 4.520 3.605 ;
        RECT  4.430 1.145 4.515 3.605 ;
        RECT  4.290 0.630 4.430 3.605 ;
        RECT  4.285 0.630 4.290 3.550 ;
        RECT  4.200 0.630 4.285 1.485 ;
        RECT  3.860 2.625 4.285 2.855 ;
        RECT  4.000 1.945 4.055 2.175 ;
        RECT  3.770 1.940 4.000 2.175 ;
        RECT  3.520 2.570 3.860 2.910 ;
        RECT  2.890 1.940 3.770 2.170 ;
        RECT  2.660 1.115 2.890 3.590 ;
        RECT  2.120 1.115 2.660 1.345 ;
        RECT  2.200 1.960 2.430 4.225 ;
        RECT  2.100 1.960 2.200 2.190 ;
        RECT  0.610 3.995 2.200 4.225 ;
        RECT  1.870 1.695 2.100 2.190 ;
        RECT  0.390 2.890 0.610 4.225 ;
        RECT  0.390 1.445 0.540 1.785 ;
        RECT  0.380 1.445 0.390 4.225 ;
        RECT  0.270 1.445 0.380 4.190 ;
        RECT  0.200 1.445 0.270 3.120 ;
        RECT  0.160 1.550 0.200 3.120 ;
    END
END DFFHQX4

MACRO DFFHQX2
    CLASS CORE ;
    FOREIGN DFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFHQXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 0.700 12.240 1.040 ;
        RECT  11.525 0.810 11.900 1.040 ;
        RECT  11.525 2.940 11.740 3.220 ;
        RECT  11.295 0.810 11.525 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 1.405 1.825 2.075 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.490 2.770 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.000 -0.400 13.200 0.400 ;
        RECT  12.660 -0.400 13.000 0.950 ;
        RECT  11.440 -0.400 12.660 0.400 ;
        RECT  11.100 -0.400 11.440 0.575 ;
        RECT  9.425 -0.400 11.100 0.400 ;
        RECT  9.195 -0.400 9.425 1.075 ;
        RECT  6.320 -0.400 9.195 0.400 ;
        RECT  5.980 -0.400 6.320 1.440 ;
        RECT  4.020 -0.400 5.980 0.400 ;
        RECT  3.680 -0.400 4.020 1.270 ;
        RECT  1.080 -0.400 3.680 0.400 ;
        RECT  0.740 -0.400 1.080 0.575 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.340 4.640 13.200 5.440 ;
        RECT  12.000 4.465 12.340 5.440 ;
        RECT  10.360 4.640 12.000 5.440 ;
        RECT  8.610 4.465 10.360 5.440 ;
        RECT  5.910 4.640 8.610 5.440 ;
        RECT  5.570 4.465 5.910 5.440 ;
        RECT  1.970 4.640 5.570 5.440 ;
        RECT  1.630 4.465 1.970 5.440 ;
        RECT  0.000 4.640 1.630 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.435 1.515 12.665 4.140 ;
        RECT  11.900 1.515 12.435 1.745 ;
        RECT  11.580 3.910 12.435 4.140 ;
        RECT  11.970 2.285 12.200 3.680 ;
        RECT  11.065 3.450 11.970 3.680 ;
        RECT  11.235 3.910 11.580 4.370 ;
        RECT  10.605 3.910 11.235 4.140 ;
        RECT  10.835 1.500 11.065 3.680 ;
        RECT  10.280 1.500 10.835 1.730 ;
        RECT  9.450 3.360 10.835 3.590 ;
        RECT  10.375 1.960 10.605 3.130 ;
        RECT  10.375 3.905 10.605 4.140 ;
        RECT  8.465 1.960 10.375 2.190 ;
        RECT  8.195 2.900 10.375 3.130 ;
        RECT  10.060 3.905 10.375 4.135 ;
        RECT  9.940 1.165 10.280 1.730 ;
        RECT  7.470 2.420 10.070 2.650 ;
        RECT  8.925 1.500 9.940 1.730 ;
        RECT  9.340 3.360 9.450 3.700 ;
        RECT  9.110 3.360 9.340 4.135 ;
        RECT  7.130 3.905 9.110 4.135 ;
        RECT  8.695 0.640 8.925 1.730 ;
        RECT  7.950 0.640 8.695 0.870 ;
        RECT  8.235 1.100 8.465 2.190 ;
        RECT  7.025 1.445 8.235 1.675 ;
        RECT  7.965 2.900 8.195 3.675 ;
        RECT  7.850 3.390 7.965 3.675 ;
        RECT  7.720 0.640 7.950 1.215 ;
        RECT  6.695 3.390 7.850 3.620 ;
        RECT  7.460 0.985 7.720 1.215 ;
        RECT  7.360 2.420 7.470 3.160 ;
        RECT  7.130 1.905 7.360 3.160 ;
        RECT  5.510 1.905 7.130 2.135 ;
        RECT  6.235 2.930 7.130 3.160 ;
        RECT  6.795 1.100 7.025 1.675 ;
        RECT  6.465 3.390 6.695 3.730 ;
        RECT  5.775 2.365 6.610 2.595 ;
        RECT  6.005 2.930 6.235 4.235 ;
        RECT  2.375 4.005 6.005 4.235 ;
        RECT  5.545 2.365 5.775 3.775 ;
        RECT  4.765 3.545 5.545 3.775 ;
        RECT  5.375 1.105 5.520 1.445 ;
        RECT  5.280 0.630 5.375 1.445 ;
        RECT  5.280 2.365 5.315 2.965 ;
        RECT  5.085 0.630 5.280 2.965 ;
        RECT  5.050 0.630 5.085 2.595 ;
        RECT  5.015 0.630 5.050 0.860 ;
        RECT  4.535 0.950 4.765 3.775 ;
        RECT  3.625 2.160 4.535 2.500 ;
        RECT  3.395 1.545 4.180 1.775 ;
        RECT  3.165 1.545 3.395 3.600 ;
        RECT  2.970 1.545 3.165 1.775 ;
        RECT  2.740 0.920 2.970 1.775 ;
        RECT  2.660 0.920 2.740 1.150 ;
        RECT  2.320 0.810 2.660 1.150 ;
        RECT  2.375 1.380 2.430 1.720 ;
        RECT  2.145 1.380 2.375 4.235 ;
        RECT  2.090 1.380 2.145 1.720 ;
        RECT  1.210 3.135 2.145 3.365 ;
        RECT  0.870 3.025 1.210 3.365 ;
        RECT  0.570 3.025 0.870 3.255 ;
        RECT  0.340 1.340 0.570 3.255 ;
        RECT  0.180 1.340 0.340 1.680 ;
    END
END DFFHQX2

MACRO DFFHQX1
    CLASS CORE ;
    FOREIGN DFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFHQXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 0.695 10.435 3.530 ;
        RECT  10.205 0.695 10.345 3.755 ;
        RECT  9.590 0.695 10.205 0.925 ;
        RECT  10.115 3.190 10.205 3.755 ;
        RECT  9.050 3.190 10.115 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 1.820 1.840 2.630 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.205 1.180 2.660 ;
        RECT  0.645 2.150 0.875 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 -0.400 10.560 0.400 ;
        RECT  8.830 -0.400 9.170 0.575 ;
        RECT  6.315 -0.400 8.830 0.400 ;
        RECT  6.085 -0.400 6.315 1.460 ;
        RECT  4.015 -0.400 6.085 0.400 ;
        RECT  3.785 -0.400 4.015 1.150 ;
        RECT  1.350 -0.400 3.785 0.400 ;
        RECT  1.010 -0.400 1.350 0.575 ;
        RECT  0.000 -0.400 1.010 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.120 4.640 10.560 5.440 ;
        RECT  9.780 4.410 10.120 5.440 ;
        RECT  8.630 4.640 9.780 5.440 ;
        RECT  8.290 4.465 8.630 5.440 ;
        RECT  5.795 4.640 8.290 5.440 ;
        RECT  5.455 4.465 5.795 5.440 ;
        RECT  1.815 4.640 5.455 5.440 ;
        RECT  1.475 4.465 1.815 5.440 ;
        RECT  0.000 4.640 1.475 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.925 1.460 9.970 1.800 ;
        RECT  9.695 1.460 9.925 2.960 ;
        RECT  9.630 1.460 9.695 1.800 ;
        RECT  8.640 2.730 9.695 2.960 ;
        RECT  9.235 2.040 9.465 2.380 ;
        RECT  9.090 4.115 9.390 4.345 ;
        RECT  9.170 2.040 9.235 2.270 ;
        RECT  8.940 1.605 9.170 2.270 ;
        RECT  8.860 4.005 9.090 4.345 ;
        RECT  7.955 1.605 8.940 1.835 ;
        RECT  8.640 4.005 8.860 4.235 ;
        RECT  8.410 2.180 8.640 4.235 ;
        RECT  8.300 2.180 8.410 2.520 ;
        RECT  6.775 0.875 8.390 1.105 ;
        RECT  7.725 1.440 7.955 4.375 ;
        RECT  7.030 4.145 7.725 4.375 ;
        RECT  7.265 1.445 7.495 3.915 ;
        RECT  7.235 1.445 7.265 1.675 ;
        RECT  6.595 3.685 7.265 3.915 ;
        RECT  7.005 1.335 7.235 1.675 ;
        RECT  6.865 2.820 7.035 3.165 ;
        RECT  6.775 1.905 6.865 3.455 ;
        RECT  6.635 0.875 6.775 3.455 ;
        RECT  6.545 0.875 6.635 2.135 ;
        RECT  6.135 3.225 6.635 3.455 ;
        RECT  6.365 3.685 6.595 4.185 ;
        RECT  5.905 1.905 6.545 2.135 ;
        RECT  6.135 2.380 6.365 2.995 ;
        RECT  5.675 2.765 6.135 2.995 ;
        RECT  5.905 3.225 6.135 4.235 ;
        RECT  5.675 1.765 5.905 2.135 ;
        RECT  2.375 4.005 5.905 4.235 ;
        RECT  5.560 1.765 5.675 1.995 ;
        RECT  5.445 2.765 5.675 3.775 ;
        RECT  5.365 1.170 5.570 1.510 ;
        RECT  4.625 3.545 5.445 3.775 ;
        RECT  5.275 0.630 5.365 1.510 ;
        RECT  5.215 0.630 5.275 1.615 ;
        RECT  5.135 0.630 5.215 3.130 ;
        RECT  5.045 1.225 5.135 3.130 ;
        RECT  4.985 1.385 5.045 3.130 ;
        RECT  4.625 0.810 4.815 1.155 ;
        RECT  4.585 0.810 4.625 3.775 ;
        RECT  4.395 0.925 4.585 3.775 ;
        RECT  3.920 2.185 4.395 2.415 ;
        RECT  3.935 1.455 4.165 1.800 ;
        RECT  3.295 1.455 3.935 1.685 ;
        RECT  3.580 2.130 3.920 2.470 ;
        RECT  3.065 0.805 3.295 3.680 ;
        RECT  2.370 0.805 3.065 1.035 ;
        RECT  2.145 1.390 2.375 4.235 ;
        RECT  1.055 3.135 2.145 3.365 ;
        RECT  0.715 3.025 1.055 3.365 ;
        RECT  0.415 1.430 0.750 1.770 ;
        RECT  0.415 3.025 0.715 3.255 ;
        RECT  0.410 1.430 0.415 3.255 ;
        RECT  0.185 1.540 0.410 3.255 ;
    END
END DFFHQX1

MACRO DFFXL
    CLASS CORE ;
    FOREIGN DFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.345 3.515 10.435 3.855 ;
        RECT  10.280 0.810 10.345 3.855 ;
        RECT  10.115 0.705 10.280 3.855 ;
        RECT  10.050 0.705 10.115 1.285 ;
        RECT  10.095 3.515 10.115 3.855 ;
        RECT  9.810 0.705 10.050 0.935 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.180 0.685 9.450 0.915 ;
        RECT  9.115 1.875 9.345 3.440 ;
        RECT  9.010 0.685 9.180 1.165 ;
        RECT  9.010 1.875 9.115 2.105 ;
        RECT  9.075 3.210 9.115 3.440 ;
        RECT  8.735 3.210 9.075 3.550 ;
        RECT  8.950 0.685 9.010 2.105 ;
        RECT  8.780 0.935 8.950 2.105 ;
        RECT  8.135 1.285 8.780 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 1.845 1.765 2.075 ;
        RECT  1.350 1.475 1.635 2.075 ;
        RECT  1.295 1.475 1.350 1.815 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.305 1.180 2.660 ;
        RECT  0.800 2.200 0.875 2.660 ;
        RECT  0.645 2.200 0.800 2.655 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.850 -0.400 11.220 0.400 ;
        RECT  10.510 -0.400 10.850 0.575 ;
        RECT  8.690 -0.400 10.510 0.400 ;
        RECT  8.350 -0.400 8.690 0.575 ;
        RECT  6.250 -0.400 8.350 0.400 ;
        RECT  5.910 -0.400 6.250 1.510 ;
        RECT  3.895 -0.400 5.910 0.400 ;
        RECT  3.665 -0.400 3.895 1.150 ;
        RECT  1.175 -0.400 3.665 0.400 ;
        RECT  0.835 -0.400 1.175 0.575 ;
        RECT  0.000 -0.400 0.835 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.735 4.640 11.220 5.440 ;
        RECT  9.395 4.410 9.735 5.440 ;
        RECT  8.275 4.640 9.395 5.440 ;
        RECT  7.935 4.465 8.275 5.440 ;
        RECT  5.795 4.640 7.935 5.440 ;
        RECT  5.455 4.465 5.795 5.440 ;
        RECT  1.380 4.640 5.455 5.440 ;
        RECT  1.040 4.410 1.380 5.440 ;
        RECT  0.000 4.640 1.040 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.580 1.415 9.810 4.180 ;
        RECT  9.240 1.415 9.580 1.645 ;
        RECT  9.095 3.950 9.580 4.180 ;
        RECT  8.865 3.950 9.095 4.350 ;
        RECT  8.645 4.005 8.865 4.350 ;
        RECT  8.310 2.670 8.795 2.900 ;
        RECT  7.850 4.005 8.645 4.235 ;
        RECT  8.080 2.260 8.310 2.900 ;
        RECT  7.530 2.260 8.080 2.490 ;
        RECT  6.775 0.670 7.930 0.900 ;
        RECT  7.620 2.745 7.850 4.235 ;
        RECT  7.240 1.270 7.530 2.490 ;
        RECT  7.190 1.270 7.240 4.150 ;
        RECT  7.115 2.260 7.190 4.150 ;
        RECT  7.010 2.260 7.115 4.260 ;
        RECT  6.775 3.920 7.010 4.260 ;
        RECT  6.665 0.670 6.775 3.260 ;
        RECT  6.545 0.670 6.665 3.615 ;
        RECT  5.665 1.740 6.545 1.970 ;
        RECT  6.435 2.920 6.545 3.615 ;
        RECT  6.270 3.385 6.435 3.615 ;
        RECT  6.205 2.200 6.310 2.690 ;
        RECT  6.040 3.385 6.270 4.235 ;
        RECT  6.080 2.200 6.205 3.135 ;
        RECT  5.975 2.460 6.080 3.135 ;
        RECT  2.790 4.005 6.040 4.235 ;
        RECT  5.800 2.905 5.975 3.135 ;
        RECT  5.570 2.905 5.800 3.775 ;
        RECT  5.590 1.740 5.665 2.325 ;
        RECT  5.435 1.740 5.590 2.510 ;
        RECT  4.660 3.545 5.570 3.775 ;
        RECT  5.245 1.170 5.450 1.510 ;
        RECT  5.360 2.095 5.435 2.510 ;
        RECT  5.175 0.630 5.245 1.510 ;
        RECT  5.130 2.780 5.235 3.120 ;
        RECT  5.130 0.630 5.175 1.610 ;
        RECT  5.015 0.630 5.130 3.120 ;
        RECT  4.945 1.225 5.015 3.120 ;
        RECT  4.900 1.380 4.945 3.120 ;
        RECT  4.895 2.780 4.900 3.120 ;
        RECT  4.660 0.810 4.695 1.150 ;
        RECT  4.465 0.810 4.660 3.775 ;
        RECT  4.430 0.920 4.465 3.775 ;
        RECT  3.865 2.455 4.430 2.685 ;
        RECT  3.375 1.785 4.200 2.015 ;
        RECT  3.525 2.400 3.865 2.740 ;
        RECT  3.250 0.795 3.375 2.015 ;
        RECT  3.020 0.795 3.250 3.680 ;
        RECT  2.250 0.795 3.020 1.025 ;
        RECT  2.560 3.250 2.790 4.235 ;
        RECT  2.315 3.250 2.560 3.480 ;
        RECT  2.085 1.390 2.315 3.480 ;
        RECT  0.540 3.250 2.085 3.480 ;
        RECT  0.380 3.140 0.540 3.480 ;
        RECT  0.380 1.065 0.520 1.405 ;
        RECT  0.200 1.065 0.380 3.480 ;
        RECT  0.180 1.065 0.200 3.370 ;
        RECT  0.150 1.120 0.180 3.370 ;
    END
END DFFXL

MACRO DFFX4
    CLASS CORE ;
    FOREIGN DFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.190 0.770 15.530 1.580 ;
        RECT  15.050 2.865 15.390 3.675 ;
        RECT  15.045 1.200 15.190 1.580 ;
        RECT  15.040 2.865 15.050 3.095 ;
        RECT  15.040 1.200 15.045 2.075 ;
        RECT  14.810 1.200 15.040 3.095 ;
        RECT  14.660 1.200 14.810 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.890 0.835 14.010 1.645 ;
        RECT  13.870 0.835 13.890 3.385 ;
        RECT  13.670 0.835 13.870 3.675 ;
        RECT  13.660 1.125 13.670 3.675 ;
        RECT  13.530 1.820 13.660 3.675 ;
        RECT  13.340 1.820 13.530 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.745 2.405 1.765 2.635 ;
        RECT  1.740 1.550 1.745 2.635 ;
        RECT  1.510 1.495 1.740 2.635 ;
        RECT  1.400 1.495 1.510 1.835 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 2.200 1.105 2.635 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.310 -0.400 16.500 0.400 ;
        RECT  15.970 -0.400 16.310 0.575 ;
        RECT  14.770 -0.400 15.970 0.400 ;
        RECT  14.430 -0.400 14.770 0.575 ;
        RECT  13.235 -0.400 14.430 0.400 ;
        RECT  13.005 -0.400 13.235 1.350 ;
        RECT  11.795 -0.400 13.005 0.400 ;
        RECT  11.565 -0.400 11.795 1.310 ;
        RECT  9.155 -0.400 11.565 0.400 ;
        RECT  8.925 -0.400 9.155 1.335 ;
        RECT  6.595 -0.400 8.925 0.400 ;
        RECT  6.365 -0.400 6.595 1.370 ;
        RECT  4.100 -0.400 6.365 0.400 ;
        RECT  3.760 -0.400 4.100 1.270 ;
        RECT  1.365 -0.400 3.760 0.400 ;
        RECT  1.025 -0.400 1.365 0.575 ;
        RECT  0.000 -0.400 1.025 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.150 4.640 16.500 5.440 ;
        RECT  15.810 4.465 16.150 5.440 ;
        RECT  14.630 4.640 15.810 5.440 ;
        RECT  14.290 4.465 14.630 5.440 ;
        RECT  13.110 4.640 14.290 5.440 ;
        RECT  12.770 4.465 13.110 5.440 ;
        RECT  11.790 4.640 12.770 5.440 ;
        RECT  11.450 4.465 11.790 5.440 ;
        RECT  9.345 4.640 11.450 5.440 ;
        RECT  9.005 4.005 9.345 5.440 ;
        RECT  6.520 4.640 9.005 5.440 ;
        RECT  6.180 4.465 6.520 5.440 ;
        RECT  3.030 4.640 6.180 5.440 ;
        RECT  2.575 4.465 3.030 5.440 ;
        RECT  1.380 4.640 2.575 5.440 ;
        RECT  1.040 4.465 1.380 5.440 ;
        RECT  0.000 4.640 1.040 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.715 2.330 15.945 4.160 ;
        RECT  15.620 2.330 15.715 2.560 ;
        RECT  13.095 3.930 15.715 4.160 ;
        RECT  15.390 2.055 15.620 2.560 ;
        RECT  12.865 2.115 13.095 4.160 ;
        RECT  12.515 2.115 12.865 2.345 ;
        RECT  12.210 3.470 12.865 3.810 ;
        RECT  12.285 1.040 12.515 2.345 ;
        RECT  11.325 2.785 12.490 3.015 ;
        RECT  11.600 2.115 12.285 2.345 ;
        RECT  11.095 0.970 11.325 3.490 ;
        RECT  10.490 0.970 11.095 1.250 ;
        RECT  10.630 3.260 11.095 3.490 ;
        RECT  10.260 1.550 10.860 1.780 ;
        RECT  10.290 3.260 10.630 4.070 ;
        RECT  10.150 0.965 10.490 1.305 ;
        RECT  8.060 3.450 10.290 3.680 ;
        RECT  10.205 1.550 10.260 2.935 ;
        RECT  10.030 1.550 10.205 2.970 ;
        RECT  9.800 1.075 10.150 1.305 ;
        RECT  9.920 2.595 10.030 2.970 ;
        RECT  9.755 2.740 9.920 2.970 ;
        RECT  9.570 1.075 9.800 1.805 ;
        RECT  9.525 2.740 9.755 3.040 ;
        RECT  8.530 1.575 9.570 1.805 ;
        RECT  8.300 2.810 9.525 3.040 ;
        RECT  9.230 2.235 9.285 2.575 ;
        RECT  8.945 2.035 9.230 2.575 ;
        RECT  7.020 2.035 8.945 2.265 ;
        RECT  8.300 1.250 8.530 1.805 ;
        RECT  7.930 1.250 8.300 1.480 ;
        RECT  8.015 2.595 8.300 3.040 ;
        RECT  7.720 3.450 8.060 4.260 ;
        RECT  7.960 2.595 8.015 3.000 ;
        RECT  6.795 2.760 7.960 3.000 ;
        RECT  7.590 1.140 7.930 1.480 ;
        RECT  6.965 2.035 7.020 2.400 ;
        RECT  6.735 1.600 6.965 2.400 ;
        RECT  6.565 2.760 6.795 4.225 ;
        RECT  6.135 1.600 6.735 1.830 ;
        RECT  6.680 2.060 6.735 2.400 ;
        RECT  6.445 2.760 6.565 2.990 ;
        RECT  3.535 3.995 6.565 4.225 ;
        RECT  6.350 2.225 6.445 2.990 ;
        RECT  6.215 2.115 6.350 2.990 ;
        RECT  6.010 2.115 6.215 2.455 ;
        RECT  5.905 0.630 6.135 1.830 ;
        RECT  5.980 3.315 6.110 3.655 ;
        RECT  5.770 2.705 5.980 3.655 ;
        RECT  4.820 0.630 5.905 0.860 ;
        RECT  5.750 2.705 5.770 3.600 ;
        RECT  5.310 2.705 5.750 2.935 ;
        RECT  5.445 1.175 5.675 1.690 ;
        RECT  5.370 1.460 5.445 1.690 ;
        RECT  5.365 1.460 5.370 2.190 ;
        RECT  5.310 1.460 5.365 2.245 ;
        RECT  5.140 1.460 5.310 2.935 ;
        RECT  4.805 3.320 5.145 3.660 ;
        RECT  5.080 1.905 5.140 2.935 ;
        RECT  5.025 1.905 5.080 2.245 ;
        RECT  4.795 0.630 4.820 1.485 ;
        RECT  4.800 3.320 4.805 3.605 ;
        RECT  4.795 2.625 4.800 3.605 ;
        RECT  4.590 0.630 4.795 3.605 ;
        RECT  4.570 1.145 4.590 3.605 ;
        RECT  4.565 1.145 4.570 3.550 ;
        RECT  4.480 1.145 4.565 1.485 ;
        RECT  4.140 2.625 4.565 2.855 ;
        RECT  4.280 1.945 4.335 2.175 ;
        RECT  4.050 1.940 4.280 2.175 ;
        RECT  3.800 2.570 4.140 2.910 ;
        RECT  3.170 1.940 4.050 2.170 ;
        RECT  3.250 3.890 3.535 4.225 ;
        RECT  2.710 3.890 3.250 4.150 ;
        RECT  2.940 0.685 3.170 3.590 ;
        RECT  2.400 0.685 2.940 0.915 ;
        RECT  2.480 2.820 2.710 4.150 ;
        RECT  2.360 2.820 2.480 3.050 ;
        RECT  1.840 3.920 2.480 4.150 ;
        RECT  2.130 1.390 2.360 3.050 ;
        RECT  1.610 3.920 1.840 4.235 ;
        RECT  0.620 4.005 1.610 4.235 ;
        RECT  0.350 2.870 0.620 4.235 ;
        RECT  0.350 0.845 0.520 1.655 ;
        RECT  0.280 0.845 0.350 4.235 ;
        RECT  0.180 0.845 0.280 3.255 ;
        RECT  0.120 1.135 0.180 3.255 ;
    END
END DFFX4

MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 1.355 12.985 3.330 ;
        RECT  12.680 1.355 12.755 1.845 ;
        RECT  12.700 3.100 12.755 3.330 ;
        RECT  12.360 3.100 12.700 3.440 ;
        RECT  12.580 1.355 12.680 1.695 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.505 0.700 11.560 1.040 ;
        RECT  11.220 0.700 11.505 1.080 ;
        RECT  10.865 0.850 11.220 1.080 ;
        RECT  11.080 2.870 11.160 3.210 ;
        RECT  10.865 2.380 11.080 3.210 ;
        RECT  10.820 0.850 10.865 3.210 ;
        RECT  10.700 0.850 10.820 2.660 ;
        RECT  10.635 0.850 10.700 2.610 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.405 1.825 2.075 ;
        RECT  1.325 1.405 1.460 1.745 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.120 1.180 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.480 -0.400 13.860 0.400 ;
        RECT  13.140 -0.400 13.480 0.575 ;
        RECT  12.360 -0.400 13.140 0.400 ;
        RECT  12.020 -0.400 12.360 0.575 ;
        RECT  10.760 -0.400 12.020 0.400 ;
        RECT  10.420 -0.400 10.760 0.575 ;
        RECT  8.800 -0.400 10.420 0.400 ;
        RECT  8.460 -0.400 8.800 1.270 ;
        RECT  6.185 -0.400 8.460 0.400 ;
        RECT  5.845 -0.400 6.185 1.445 ;
        RECT  4.020 -0.400 5.845 0.400 ;
        RECT  3.680 -0.400 4.020 1.270 ;
        RECT  1.100 -0.400 3.680 0.400 ;
        RECT  0.760 -0.400 1.100 0.575 ;
        RECT  0.000 -0.400 0.760 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.260 4.640 13.860 5.440 ;
        RECT  12.920 4.465 13.260 5.440 ;
        RECT  11.920 4.640 12.920 5.440 ;
        RECT  11.580 4.465 11.920 5.440 ;
        RECT  9.940 4.640 11.580 5.440 ;
        RECT  8.190 4.465 9.940 5.440 ;
        RECT  5.890 4.640 8.190 5.440 ;
        RECT  5.550 4.465 5.890 5.440 ;
        RECT  4.530 4.640 5.550 5.440 ;
        RECT  4.190 4.465 4.530 5.440 ;
        RECT  1.450 4.640 4.190 5.440 ;
        RECT  1.110 4.410 1.450 5.440 ;
        RECT  0.000 4.640 1.110 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.435 4.020 12.490 4.360 ;
        RECT  12.150 3.995 12.435 4.360 ;
        RECT  12.125 3.995 12.150 4.225 ;
        RECT  11.895 1.545 12.125 4.225 ;
        RECT  11.220 1.545 11.895 1.775 ;
        RECT  11.160 3.995 11.895 4.225 ;
        RECT  11.435 2.285 11.665 3.670 ;
        RECT  9.975 3.440 11.435 3.670 ;
        RECT  11.050 3.995 11.160 4.370 ;
        RECT  10.820 3.900 11.050 4.370 ;
        RECT  9.640 3.900 10.820 4.130 ;
        RECT  9.745 1.775 9.975 3.670 ;
        RECT  9.600 1.775 9.745 2.005 ;
        RECT  9.030 3.360 9.745 3.670 ;
        RECT  9.370 1.155 9.600 2.005 ;
        RECT  9.110 2.350 9.450 2.690 ;
        RECT  9.260 1.155 9.370 1.795 ;
        RECT  8.130 1.565 9.260 1.795 ;
        RECT  8.195 2.405 9.110 2.635 ;
        RECT  8.920 3.360 9.030 3.700 ;
        RECT  8.690 3.360 8.920 3.960 ;
        RECT  7.155 3.730 8.690 3.960 ;
        RECT  7.965 2.405 8.195 3.160 ;
        RECT  7.900 1.160 8.130 1.795 ;
        RECT  7.300 2.930 7.965 3.160 ;
        RECT  7.520 1.160 7.900 1.390 ;
        RECT  7.180 1.050 7.520 1.390 ;
        RECT  7.210 2.820 7.300 3.160 ;
        RECT  6.980 1.785 7.210 3.160 ;
        RECT  6.925 3.440 7.155 4.275 ;
        RECT  5.530 1.785 6.980 2.015 ;
        RECT  6.960 2.820 6.980 3.160 ;
        RECT  6.330 2.930 6.960 3.160 ;
        RECT  5.860 2.245 6.610 2.475 ;
        RECT  6.100 2.930 6.330 4.235 ;
        RECT  3.595 4.005 6.100 4.235 ;
        RECT  5.630 2.245 5.860 3.775 ;
        RECT  4.695 3.545 5.630 3.775 ;
        RECT  5.295 1.105 5.445 1.445 ;
        RECT  5.295 2.625 5.330 2.965 ;
        RECT  5.065 0.630 5.295 2.965 ;
        RECT  4.935 0.630 5.065 0.860 ;
        RECT  4.990 2.625 5.065 2.965 ;
        RECT  4.685 2.270 4.695 3.775 ;
        RECT  4.465 0.950 4.685 3.775 ;
        RECT  4.455 0.950 4.465 2.510 ;
        RECT  3.585 2.170 4.455 2.510 ;
        RECT  3.355 1.555 4.180 1.785 ;
        RECT  3.365 3.890 3.595 4.235 ;
        RECT  3.310 3.890 3.365 4.225 ;
        RECT  3.125 1.545 3.355 3.600 ;
        RECT  3.300 3.890 3.310 4.150 ;
        RECT  2.895 3.890 3.300 4.120 ;
        RECT  2.970 1.545 3.125 1.785 ;
        RECT  2.740 0.920 2.970 1.785 ;
        RECT  2.665 2.820 2.895 4.120 ;
        RECT  2.660 0.920 2.740 1.150 ;
        RECT  2.375 2.820 2.665 3.050 ;
        RECT  1.980 3.890 2.665 4.120 ;
        RECT  2.320 0.810 2.660 1.150 ;
        RECT  2.375 1.380 2.430 1.720 ;
        RECT  2.145 1.380 2.375 3.050 ;
        RECT  2.090 1.380 2.145 1.720 ;
        RECT  1.750 3.605 1.980 4.120 ;
        RECT  1.310 3.605 1.750 3.835 ;
        RECT  0.910 3.020 1.310 3.835 ;
        RECT  0.570 3.080 0.910 3.310 ;
        RECT  0.340 1.340 0.570 3.310 ;
        RECT  0.180 1.340 0.340 1.680 ;
    END
END DFFX2

MACRO DFFX1
    CLASS CORE ;
    FOREIGN DFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 1.190 11.040 3.880 ;
        RECT  10.600 3.540 10.700 3.880 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 0.865 10.345 3.420 ;
        RECT  9.830 0.865 10.115 1.095 ;
        RECT  9.230 3.190 10.115 3.420 ;
        RECT  9.300 0.695 9.830 1.095 ;
        RECT  8.890 3.190 9.230 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 1.845 1.765 2.075 ;
        RECT  1.410 1.405 1.690 2.075 ;
        RECT  1.290 1.405 1.410 1.745 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER METAL1 ;
        RECT  0.940 2.205 1.180 2.660 ;
        RECT  0.710 2.150 0.940 2.660 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.460 -0.400 11.220 0.400 ;
        RECT  10.120 -0.400 10.460 0.575 ;
        RECT  8.880 -0.400 10.120 0.400 ;
        RECT  8.540 -0.400 8.880 0.575 ;
        RECT  6.440 -0.400 8.540 0.400 ;
        RECT  6.100 -0.400 6.440 1.460 ;
        RECT  4.015 -0.400 6.100 0.400 ;
        RECT  3.785 -0.400 4.015 1.150 ;
        RECT  1.225 -0.400 3.785 0.400 ;
        RECT  0.885 -0.400 1.225 0.575 ;
        RECT  0.000 -0.400 0.885 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.180 4.640 11.220 5.440 ;
        RECT  9.840 4.410 10.180 5.440 ;
        RECT  8.470 4.640 9.840 5.440 ;
        RECT  8.130 4.465 8.470 5.440 ;
        RECT  5.795 4.640 8.130 5.440 ;
        RECT  5.455 4.465 5.795 5.440 ;
        RECT  1.550 4.640 5.455 5.440 ;
        RECT  1.210 4.465 1.550 5.440 ;
        RECT  0.000 4.640 1.210 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.680 1.600 9.870 2.765 ;
        RECT  9.640 1.490 9.680 2.765 ;
        RECT  9.340 1.490 9.640 1.830 ;
        RECT  8.400 2.535 9.640 2.765 ;
        RECT  8.880 2.075 9.255 2.305 ;
        RECT  9.110 4.140 9.230 4.370 ;
        RECT  8.880 3.970 9.110 4.370 ;
        RECT  8.650 1.440 8.880 2.305 ;
        RECT  8.400 3.970 8.880 4.200 ;
        RECT  7.550 1.440 8.650 1.835 ;
        RECT  8.350 2.535 8.400 4.200 ;
        RECT  8.170 2.180 8.350 4.200 ;
        RECT  8.120 2.180 8.170 2.765 ;
        RECT  8.010 2.180 8.120 2.520 ;
        RECT  6.940 0.875 8.100 1.105 ;
        RECT  7.320 1.440 7.550 4.285 ;
        RECT  6.870 4.055 7.320 4.285 ;
        RECT  6.940 2.820 7.090 3.160 ;
        RECT  6.865 0.875 6.940 3.160 ;
        RECT  6.710 0.875 6.865 3.615 ;
        RECT  6.635 1.765 6.710 3.615 ;
        RECT  5.560 1.765 6.635 1.995 ;
        RECT  6.270 3.385 6.635 3.615 ;
        RECT  6.135 2.380 6.365 3.135 ;
        RECT  6.040 3.385 6.270 4.235 ;
        RECT  5.800 2.905 6.135 3.135 ;
        RECT  3.535 4.005 6.040 4.235 ;
        RECT  5.570 2.905 5.800 3.775 ;
        RECT  5.405 1.170 5.610 1.510 ;
        RECT  4.760 3.545 5.570 3.775 ;
        RECT  5.315 0.630 5.405 1.510 ;
        RECT  5.315 2.790 5.330 3.130 ;
        RECT  5.085 0.630 5.315 3.130 ;
        RECT  4.990 2.790 5.085 3.130 ;
        RECT  4.760 0.810 4.815 2.470 ;
        RECT  4.585 0.810 4.760 3.775 ;
        RECT  4.490 2.130 4.585 3.775 ;
        RECT  3.580 2.130 4.490 2.470 ;
        RECT  3.375 1.515 4.355 1.745 ;
        RECT  2.835 3.995 3.535 4.235 ;
        RECT  3.295 0.805 3.375 1.745 ;
        RECT  3.065 0.805 3.295 3.680 ;
        RECT  2.370 0.805 3.065 1.035 ;
        RECT  2.605 2.820 2.835 4.235 ;
        RECT  2.375 2.820 2.605 3.050 ;
        RECT  0.785 3.605 2.605 3.835 ;
        RECT  2.145 1.390 2.375 3.050 ;
        RECT  0.445 3.020 0.785 3.835 ;
        RECT  0.445 1.430 0.520 1.770 ;
        RECT  0.365 1.430 0.445 3.835 ;
        RECT  0.215 1.430 0.365 3.310 ;
        RECT  0.180 1.430 0.215 1.770 ;
    END
END DFFX1

MACRO CLKINVXL
    CLASS CORE ;
    FOREIGN CLKINVXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 1.820 1.830 3.220 ;
        RECT  1.255 1.350 1.485 3.885 ;
        RECT  1.120 1.350 1.255 1.850 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.190 2.380 0.925 2.810 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 -0.400 1.980 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.890 4.640 1.980 5.440 ;
        RECT  0.525 4.395 0.890 5.440 ;
        RECT  0.000 4.640 0.525 5.440 ;
        END
    END VDD
END CLKINVXL

MACRO CLKINVX8
    CLASS CORE ;
    FOREIGN CLKINVX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 1.820 3.745 3.220 ;
        RECT  3.085 1.510 3.160 3.220 ;
        RECT  2.880 1.510 3.085 3.275 ;
        RECT  2.195 1.235 2.880 3.410 ;
        RECT  2.120 1.235 2.195 1.820 ;
        RECT  0.780 2.930 2.195 3.410 ;
        RECT  0.870 1.235 2.120 1.715 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.045 1.355 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 -0.400 3.960 0.400 ;
        RECT  1.665 -0.400 2.005 0.980 ;
        RECT  0.560 -0.400 1.665 0.400 ;
        RECT  0.220 -0.400 0.560 0.575 ;
        RECT  0.000 -0.400 0.220 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 4.640 3.960 5.440 ;
        RECT  2.980 3.790 3.320 5.440 ;
        RECT  1.915 4.640 2.980 5.440 ;
        RECT  1.575 3.790 1.915 5.440 ;
        RECT  0.520 4.640 1.575 5.440 ;
        RECT  0.180 3.790 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END CLKINVX8

MACRO CLKINVX4
    CLASS CORE ;
    FOREIGN CLKINVX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.290 1.840 3.780 ;
        RECT  1.080 1.290 1.460 1.670 ;
        RECT  1.440 2.965 1.460 3.780 ;
        RECT  1.100 2.965 1.440 4.205 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.020 0.950 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 -0.400 2.640 0.400 ;
        RECT  2.100 -0.400 2.440 0.575 ;
        RECT  0.680 -0.400 2.100 0.400 ;
        RECT  0.340 -0.400 0.680 0.575 ;
        RECT  0.000 -0.400 0.340 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 4.640 2.640 5.440 ;
        RECT  1.860 4.465 2.200 5.440 ;
        RECT  0.680 4.640 1.860 5.440 ;
        RECT  0.340 4.465 0.680 5.440 ;
        RECT  0.000 4.640 0.340 5.440 ;
        END
    END VDD
END CLKINVX4

MACRO CLKINVX3
    CLASS CORE ;
    FOREIGN CLKINVX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.025 2.630 1.180 3.780 ;
        RECT  0.795 1.435 1.025 3.780 ;
        RECT  0.735 2.635 0.795 3.780 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.535 2.440 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 -0.400 1.980 0.400 ;
        RECT  1.300 -0.400 1.640 0.575 ;
        RECT  0.000 -0.400 1.300 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 4.640 1.980 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
END CLKINVX3

MACRO CLKINVX2
    CLASS CORE ;
    FOREIGN CLKINVX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 1.200 1.550 3.305 ;
        RECT  1.155 1.200 1.320 1.540 ;
        RECT  0.740 2.940 1.320 3.305 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 1.085 2.410 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 -0.400 1.980 0.400 ;
        RECT  0.385 -0.400 0.725 1.540 ;
        RECT  0.000 -0.400 0.385 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.450 4.640 1.980 5.440 ;
        RECT  1.070 4.395 1.450 5.440 ;
        RECT  0.000 4.640 1.070 5.440 ;
        END
    END VDD
END CLKINVX2

MACRO CLKINVX20
    CLASS CORE ;
    FOREIGN CLKINVX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.265 2.925 18.890 3.735 ;
        RECT  16.715 1.200 18.265 3.780 ;
        RECT  15.115 1.200 16.715 1.880 ;
        RECT  16.055 2.990 16.715 3.670 ;
        RECT  15.490 2.925 16.055 3.735 ;
        RECT  14.735 2.990 15.490 3.670 ;
        RECT  13.640 1.195 15.115 1.880 ;
        RECT  14.120 2.925 14.735 3.735 ;
        RECT  13.055 2.990 14.120 3.670 ;
        RECT  10.660 1.200 13.640 1.880 ;
        RECT  12.715 2.925 13.055 3.735 ;
        RECT  11.620 2.990 12.715 3.670 ;
        RECT  11.005 2.925 11.620 3.735 ;
        RECT  10.200 2.990 11.005 3.670 ;
        RECT  10.320 1.195 10.660 1.880 ;
        RECT  8.900 1.195 10.320 1.875 ;
        RECT  9.685 2.925 10.200 3.735 ;
        RECT  8.795 2.990 9.685 3.670 ;
        RECT  8.365 2.925 8.795 3.735 ;
        RECT  7.475 2.990 8.365 3.670 ;
        RECT  7.010 2.925 7.475 3.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.715 2.100 1.180 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.780 -0.400 19.140 0.400 ;
        RECT  15.440 -0.400 15.780 0.960 ;
        RECT  14.395 -0.400 15.440 0.400 ;
        RECT  14.055 -0.400 14.395 0.960 ;
        RECT  12.975 -0.400 14.055 0.400 ;
        RECT  12.635 -0.400 12.975 0.960 ;
        RECT  11.545 -0.400 12.635 0.400 ;
        RECT  11.205 -0.400 11.545 0.960 ;
        RECT  10.125 -0.400 11.205 0.400 ;
        RECT  9.785 -0.400 10.125 0.960 ;
        RECT  8.705 -0.400 9.785 0.400 ;
        RECT  8.365 -0.400 8.705 0.960 ;
        RECT  5.185 -0.400 8.365 0.400 ;
        RECT  4.845 -0.400 5.185 0.945 ;
        RECT  3.640 -0.400 4.845 0.400 ;
        RECT  3.300 -0.400 3.640 0.945 ;
        RECT  2.215 -0.400 3.300 0.400 ;
        RECT  1.875 -0.400 2.215 1.000 ;
        RECT  0.000 -0.400 1.875 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.015 4.640 19.140 5.440 ;
        RECT  17.675 4.120 18.015 5.440 ;
        RECT  16.590 4.640 17.675 5.440 ;
        RECT  16.250 4.120 16.590 5.440 ;
        RECT  15.170 4.640 16.250 5.440 ;
        RECT  14.830 4.120 15.170 5.440 ;
        RECT  13.745 4.640 14.830 5.440 ;
        RECT  13.405 4.120 13.745 5.440 ;
        RECT  12.335 4.640 13.405 5.440 ;
        RECT  11.995 4.120 12.335 5.440 ;
        RECT  10.915 4.640 11.995 5.440 ;
        RECT  10.575 4.065 10.915 5.440 ;
        RECT  9.480 4.640 10.575 5.440 ;
        RECT  9.140 4.065 9.480 5.440 ;
        RECT  8.060 4.640 9.140 5.440 ;
        RECT  7.720 4.065 8.060 5.440 ;
        RECT  6.640 4.640 7.720 5.440 ;
        RECT  6.300 4.075 6.640 5.440 ;
        RECT  5.070 4.640 6.300 5.440 ;
        RECT  4.730 4.060 5.070 5.440 ;
        RECT  3.635 4.640 4.730 5.440 ;
        RECT  3.295 4.060 3.635 5.440 ;
        RECT  2.165 4.640 3.295 5.440 ;
        RECT  1.825 4.090 2.165 5.440 ;
        RECT  0.805 4.640 1.825 5.440 ;
        RECT  0.465 3.050 0.805 5.440 ;
        RECT  0.000 4.640 0.465 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 2.120 16.205 2.690 ;
        RECT  5.805 1.180 6.345 3.450 ;
        RECT  5.700 1.180 5.805 3.675 ;
        RECT  2.590 1.180 5.700 1.825 ;
        RECT  5.465 2.805 5.700 3.675 ;
        RECT  4.345 2.805 5.465 3.450 ;
        RECT  2.365 2.100 5.055 2.440 ;
        RECT  4.005 2.805 4.345 3.735 ;
        RECT  2.925 2.805 4.005 3.450 ;
        RECT  2.590 2.805 2.925 3.735 ;
        RECT  2.585 2.925 2.590 3.735 ;
        RECT  1.640 2.155 2.365 2.385 ;
        RECT  1.410 1.440 1.640 3.315 ;
        RECT  1.225 1.440 1.410 1.780 ;
        RECT  1.235 2.975 1.410 3.315 ;
    END
END CLKINVX20

MACRO CLKINVX1
    CLASS CORE ;
    FOREIGN CLKINVX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 1.820 1.830 3.220 ;
        RECT  1.255 1.350 1.485 3.885 ;
        RECT  1.040 1.350 1.255 1.855 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.190 2.380 0.925 2.810 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 -0.400 1.980 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.890 4.640 1.980 5.440 ;
        RECT  0.525 4.395 0.890 5.440 ;
        RECT  0.000 4.640 0.525 5.440 ;
        END
    END VDD
END CLKINVX1

MACRO CLKINVX16
    CLASS CORE ;
    FOREIGN CLKINVX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.735 1.200 16.285 3.840 ;
        RECT  12.990 1.200 14.735 1.880 ;
        RECT  14.195 2.990 14.735 3.670 ;
        RECT  13.645 2.925 14.195 3.735 ;
        RECT  12.790 2.990 13.645 3.670 ;
        RECT  11.705 1.195 12.990 1.880 ;
        RECT  12.325 2.925 12.790 3.735 ;
        RECT  11.435 2.990 12.325 3.670 ;
        RECT  8.195 1.200 11.705 1.880 ;
        RECT  11.005 2.925 11.435 3.735 ;
        RECT  10.115 2.990 11.005 3.670 ;
        RECT  9.595 2.925 10.115 3.735 ;
        RECT  8.795 2.990 9.595 3.670 ;
        RECT  8.165 2.925 8.795 3.735 ;
        RECT  7.085 2.990 8.165 3.670 ;
        RECT  6.745 2.925 7.085 3.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.715 2.100 1.180 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.655 -0.400 16.500 0.400 ;
        RECT  13.315 -0.400 13.655 0.960 ;
        RECT  12.270 -0.400 13.315 0.400 ;
        RECT  11.930 -0.400 12.270 0.960 ;
        RECT  10.850 -0.400 11.930 0.400 ;
        RECT  10.510 -0.400 10.850 0.960 ;
        RECT  9.420 -0.400 10.510 0.400 ;
        RECT  9.080 -0.400 9.420 0.960 ;
        RECT  8.000 -0.400 9.080 0.400 ;
        RECT  7.660 -0.400 8.000 0.960 ;
        RECT  3.640 -0.400 7.660 0.400 ;
        RECT  3.300 -0.400 3.640 1.020 ;
        RECT  2.215 -0.400 3.300 0.400 ;
        RECT  1.875 -0.400 2.215 1.000 ;
        RECT  0.000 -0.400 1.875 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.240 4.640 16.500 5.440 ;
        RECT  15.900 4.120 16.240 5.440 ;
        RECT  14.905 4.640 15.900 5.440 ;
        RECT  14.565 4.120 14.905 5.440 ;
        RECT  13.480 4.640 14.565 5.440 ;
        RECT  13.140 4.120 13.480 5.440 ;
        RECT  12.070 4.640 13.140 5.440 ;
        RECT  11.730 4.120 12.070 5.440 ;
        RECT  10.650 4.640 11.730 5.440 ;
        RECT  10.310 4.065 10.650 5.440 ;
        RECT  9.215 4.640 10.310 5.440 ;
        RECT  8.875 4.065 9.215 5.440 ;
        RECT  7.795 4.640 8.875 5.440 ;
        RECT  7.455 4.065 7.795 5.440 ;
        RECT  6.375 4.640 7.455 5.440 ;
        RECT  6.035 4.075 6.375 5.440 ;
        RECT  5.070 4.640 6.035 5.440 ;
        RECT  4.730 4.060 5.070 5.440 ;
        RECT  3.635 4.640 4.730 5.440 ;
        RECT  3.295 4.060 3.635 5.440 ;
        RECT  2.165 4.640 3.295 5.440 ;
        RECT  1.825 4.090 2.165 5.440 ;
        RECT  0.805 4.640 1.825 5.440 ;
        RECT  0.465 3.050 0.805 5.440 ;
        RECT  0.000 4.640 0.465 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.440 2.190 14.300 2.530 ;
        RECT  6.020 2.210 6.440 2.510 ;
        RECT  5.340 1.340 6.020 3.390 ;
        RECT  2.585 1.340 5.340 1.870 ;
        RECT  4.345 2.700 5.340 3.390 ;
        RECT  2.275 2.100 4.965 2.440 ;
        RECT  4.005 2.700 4.345 3.735 ;
        RECT  2.925 2.700 4.005 3.390 ;
        RECT  2.585 2.700 2.925 3.735 ;
        RECT  1.640 2.155 2.275 2.385 ;
        RECT  1.410 1.440 1.640 3.315 ;
        RECT  1.225 1.440 1.410 1.780 ;
        RECT  1.235 2.975 1.410 3.315 ;
    END
END CLKINVX16

MACRO CLKINVX12
    CLASS CORE ;
    FOREIGN CLKINVX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.775 1.195 12.325 3.780 ;
        RECT  7.020 1.195 10.775 1.875 ;
        RECT  10.115 2.990 10.775 3.670 ;
        RECT  9.685 2.925 10.115 3.735 ;
        RECT  8.795 2.990 9.685 3.670 ;
        RECT  8.295 2.925 8.795 3.735 ;
        RECT  7.475 2.990 8.295 3.670 ;
        RECT  6.865 2.925 7.475 3.735 ;
        RECT  5.785 2.990 6.865 3.670 ;
        RECT  5.445 2.925 5.785 3.735 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 2.100 1.105 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.925 -0.400 12.540 0.400 ;
        RECT  10.585 -0.400 10.925 0.960 ;
        RECT  9.495 -0.400 10.585 0.400 ;
        RECT  9.155 -0.400 9.495 0.960 ;
        RECT  8.075 -0.400 9.155 0.400 ;
        RECT  7.735 -0.400 8.075 0.960 ;
        RECT  6.680 -0.400 7.735 0.400 ;
        RECT  6.340 -0.400 6.680 0.960 ;
        RECT  3.550 -0.400 6.340 0.400 ;
        RECT  3.210 -0.400 3.550 1.020 ;
        RECT  0.695 -0.400 3.210 0.400 ;
        RECT  0.355 -0.400 0.695 1.685 ;
        RECT  0.000 -0.400 0.355 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.200 4.640 12.540 5.440 ;
        RECT  11.860 4.120 12.200 5.440 ;
        RECT  10.765 4.640 11.860 5.440 ;
        RECT  10.425 4.120 10.765 5.440 ;
        RECT  9.350 4.640 10.425 5.440 ;
        RECT  9.010 4.065 9.350 5.440 ;
        RECT  7.915 4.640 9.010 5.440 ;
        RECT  7.575 4.065 7.915 5.440 ;
        RECT  6.495 4.640 7.575 5.440 ;
        RECT  6.155 4.065 6.495 5.440 ;
        RECT  5.090 4.640 6.155 5.440 ;
        RECT  4.750 4.075 5.090 5.440 ;
        RECT  3.545 4.640 4.750 5.440 ;
        RECT  3.205 4.060 3.545 5.440 ;
        RECT  2.075 4.640 3.205 5.440 ;
        RECT  1.735 4.090 2.075 5.440 ;
        RECT  0.675 4.640 1.735 5.440 ;
        RECT  0.335 2.890 0.675 5.440 ;
        RECT  0.000 4.640 0.335 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.100 2.190 10.410 2.530 ;
        RECT  4.800 1.420 5.100 3.245 ;
        RECT  4.250 1.420 4.800 1.720 ;
        RECT  4.255 2.945 4.800 3.245 ;
        RECT  2.060 2.100 4.280 2.440 ;
        RECT  3.915 2.925 4.255 3.735 ;
        RECT  2.500 1.420 4.250 1.760 ;
        RECT  2.835 2.925 3.915 3.265 ;
        RECT  2.495 2.925 2.835 3.735 ;
        RECT  1.640 2.155 2.060 2.385 ;
        RECT  1.485 1.305 1.640 3.260 ;
        RECT  1.415 1.305 1.485 3.315 ;
        RECT  1.410 1.250 1.415 3.315 ;
        RECT  1.075 1.250 1.410 1.590 ;
        RECT  1.145 2.975 1.410 3.315 ;
    END
END CLKINVX12

MACRO CLKBUFXL
    CLASS CORE ;
    FOREIGN CLKBUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 1.220 2.425 2.990 ;
        RECT  1.920 1.220 2.195 1.450 ;
        RECT  2.120 2.635 2.195 2.990 ;
        RECT  1.880 2.760 2.120 2.990 ;
        RECT  1.580 1.110 1.920 1.450 ;
        RECT  1.540 2.760 1.880 3.100 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.810 2.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 4.640 2.640 5.440 ;
        RECT  0.880 4.465 1.220 5.440 ;
        RECT  0.000 4.640 0.880 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.270 1.820 1.520 2.160 ;
        RECT  1.040 1.220 1.270 2.990 ;
        RECT  0.520 1.220 1.040 1.450 ;
        RECT  0.520 2.760 1.040 2.990 ;
        RECT  0.180 1.110 0.520 1.450 ;
        RECT  0.180 2.760 0.520 3.100 ;
    END
END CLKBUFXL

MACRO CLKBUFX8
    CLASS CORE ;
    FOREIGN CLKBUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.820 4.405 3.220 ;
        RECT  2.855 1.350 4.000 3.220 ;
        RECT  2.780 1.350 2.855 1.850 ;
        RECT  2.780 2.625 2.855 3.180 ;
        RECT  2.260 1.350 2.780 1.690 ;
        RECT  2.180 2.840 2.780 3.180 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 1.990 1.390 2.330 ;
        RECT  0.875 1.845 1.105 2.330 ;
        RECT  0.570 1.990 0.875 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 -0.400 4.620 0.400 ;
        RECT  2.900 -0.400 3.240 0.965 ;
        RECT  1.960 -0.400 2.900 0.400 ;
        RECT  1.620 -0.400 1.960 0.965 ;
        RECT  0.000 -0.400 1.620 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 4.640 4.620 5.440 ;
        RECT  4.100 3.620 4.440 5.440 ;
        RECT  3.160 4.640 4.100 5.440 ;
        RECT  2.820 3.620 3.160 5.440 ;
        RECT  1.840 4.640 2.820 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.520 4.640 1.500 5.440 ;
        RECT  0.180 3.480 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.950 2.180 2.550 2.520 ;
        RECT  1.720 1.260 1.950 2.990 ;
        RECT  1.240 1.260 1.720 1.490 ;
        RECT  1.160 2.760 1.720 2.990 ;
        RECT  0.900 1.150 1.240 1.490 ;
        RECT  0.820 2.760 1.160 3.100 ;
    END
END CLKBUFX8

MACRO CLKBUFX4
    CLASS CORE ;
    FOREIGN CLKBUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 1.260 2.500 2.660 ;
        RECT  2.120 1.260 2.350 3.000 ;
        RECT  1.700 1.390 2.120 1.730 ;
        RECT  2.040 2.770 2.120 3.000 ;
        RECT  1.700 2.770 2.040 3.110 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.810 2.395 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 -0.400 3.300 0.400 ;
        RECT  2.460 -0.400 2.800 0.575 ;
        RECT  1.180 -0.400 2.460 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 4.640 3.300 5.440 ;
        RECT  2.460 4.465 2.800 5.440 ;
        RECT  1.280 4.640 2.460 5.440 ;
        RECT  1.225 4.465 1.280 5.440 ;
        RECT  0.995 4.410 1.225 5.440 ;
        RECT  0.940 4.465 0.995 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.270 2.060 1.890 2.400 ;
        RECT  1.040 1.360 1.270 2.970 ;
        RECT  0.520 1.360 1.040 1.590 ;
        RECT  0.520 2.740 1.040 2.970 ;
        RECT  0.180 1.250 0.520 1.590 ;
        RECT  0.180 2.740 0.520 3.080 ;
    END
END CLKBUFX4

MACRO CLKBUFX3
    CLASS CORE ;
    FOREIGN CLKBUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.205 1.880 1.545 ;
        RECT  1.770 1.820 1.840 3.160 ;
        RECT  1.540 1.205 1.770 3.160 ;
        RECT  1.500 1.820 1.540 3.160 ;
        RECT  1.460 1.820 1.500 2.660 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.555 2.360 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 -0.400 2.640 0.400 ;
        RECT  2.120 -0.400 2.460 0.575 ;
        RECT  1.180 -0.400 2.120 0.400 ;
        RECT  0.840 -0.400 1.180 0.575 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 4.640 2.640 5.440 ;
        RECT  2.120 4.465 2.460 5.440 ;
        RECT  1.195 4.640 2.120 5.440 ;
        RECT  0.810 4.465 1.195 5.440 ;
        RECT  0.000 4.640 0.810 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.115 1.975 1.225 2.315 ;
        RECT  0.885 1.135 1.115 3.155 ;
        RECT  0.520 1.135 0.885 1.365 ;
        RECT  0.520 2.925 0.885 3.155 ;
        RECT  0.180 1.025 0.520 1.365 ;
        RECT  0.180 2.925 0.520 3.265 ;
    END
END CLKBUFX3

MACRO CLKBUFX2
    CLASS CORE ;
    FOREIGN CLKBUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 1.265 2.425 2.980 ;
        RECT  2.195 1.155 2.200 2.980 ;
        RECT  1.640 1.155 2.195 1.495 ;
        RECT  2.120 2.635 2.195 3.090 ;
        RECT  1.600 2.750 2.120 3.090 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.900 2.260 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 -0.400 2.640 0.400 ;
        RECT  0.880 -0.400 1.220 0.575 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 2.640 5.440 ;
        RECT  1.125 4.465 1.180 5.440 ;
        RECT  0.895 4.410 1.125 5.440 ;
        RECT  0.840 4.465 0.895 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.370 2.060 1.620 2.400 ;
        RECT  1.140 1.265 1.370 2.980 ;
        RECT  0.620 1.265 1.140 1.495 ;
        RECT  0.620 2.750 1.140 2.980 ;
        RECT  0.280 1.155 0.620 1.495 ;
        RECT  0.280 2.750 0.620 3.090 ;
    END
END CLKBUFX2

MACRO CLKBUFX20
    CLASS CORE ;
    FOREIGN CLKBUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.760 1.200 14.965 3.840 ;
        RECT  13.415 1.125 14.760 3.840 ;
        RECT  4.700 1.125 13.415 1.925 ;
        RECT  13.340 2.660 13.415 3.525 ;
        RECT  4.660 2.725 13.340 3.525 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 1.990 3.740 2.330 ;
        RECT  2.855 1.845 3.085 2.330 ;
        RECT  0.580 1.990 2.855 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.800 -0.400 15.840 0.400 ;
        RECT  10.460 -0.400 10.800 0.895 ;
        RECT  9.520 -0.400 10.460 0.400 ;
        RECT  9.180 -0.400 9.520 0.895 ;
        RECT  8.240 -0.400 9.180 0.400 ;
        RECT  7.900 -0.400 8.240 0.895 ;
        RECT  6.960 -0.400 7.900 0.400 ;
        RECT  6.620 -0.400 6.960 0.895 ;
        RECT  5.680 -0.400 6.620 0.400 ;
        RECT  5.340 -0.400 5.680 0.895 ;
        RECT  4.400 -0.400 5.340 0.400 ;
        RECT  4.060 -0.400 4.400 0.960 ;
        RECT  2.960 -0.400 4.060 0.400 ;
        RECT  2.620 -0.400 2.960 0.960 ;
        RECT  1.520 -0.400 2.620 0.400 ;
        RECT  1.180 -0.400 1.520 0.960 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.640 4.640 15.840 5.440 ;
        RECT  14.585 4.465 14.640 5.440 ;
        RECT  14.355 4.410 14.585 5.440 ;
        RECT  14.300 4.465 14.355 5.440 ;
        RECT  13.320 4.640 14.300 5.440 ;
        RECT  12.980 4.090 13.320 5.440 ;
        RECT  12.040 4.640 12.980 5.440 ;
        RECT  11.700 4.090 12.040 5.440 ;
        RECT  10.760 4.640 11.700 5.440 ;
        RECT  10.420 4.090 10.760 5.440 ;
        RECT  9.480 4.640 10.420 5.440 ;
        RECT  9.140 4.090 9.480 5.440 ;
        RECT  8.200 4.640 9.140 5.440 ;
        RECT  7.860 4.090 8.200 5.440 ;
        RECT  6.920 4.640 7.860 5.440 ;
        RECT  6.580 4.020 6.920 5.440 ;
        RECT  5.640 4.640 6.580 5.440 ;
        RECT  5.300 4.020 5.640 5.440 ;
        RECT  4.360 4.640 5.300 5.440 ;
        RECT  4.020 3.945 4.360 5.440 ;
        RECT  3.080 4.640 4.020 5.440 ;
        RECT  2.740 3.945 3.080 5.440 ;
        RECT  1.800 4.640 2.740 5.440 ;
        RECT  1.460 3.945 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.945 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.420 2.155 12.920 2.495 ;
        RECT  4.080 1.190 4.420 3.180 ;
        RECT  1.900 1.190 4.080 1.530 ;
        RECT  0.820 2.840 4.080 3.180 ;
    END
END CLKBUFX20

MACRO CLKBUFX1
    CLASS CORE ;
    FOREIGN CLKBUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 1.220 2.425 3.050 ;
        RECT  1.920 1.220 2.195 1.450 ;
        RECT  2.120 2.635 2.195 3.050 ;
        RECT  1.840 2.820 2.120 3.050 ;
        RECT  1.580 1.110 1.920 1.450 ;
        RECT  1.500 2.820 1.840 3.160 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.810 2.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 2.640 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.270 2.060 1.520 2.400 ;
        RECT  1.040 1.220 1.270 2.990 ;
        RECT  0.520 1.220 1.040 1.450 ;
        RECT  0.520 2.760 1.040 2.990 ;
        RECT  0.180 1.110 0.520 1.450 ;
        RECT  0.180 2.760 0.520 3.100 ;
    END
END CLKBUFX1

MACRO CLKBUFX16
    CLASS CORE ;
    FOREIGN CLKBUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.120 1.200 12.325 3.840 ;
        RECT  10.775 1.125 12.120 3.840 ;
        RECT  4.060 1.125 10.775 1.925 ;
        RECT  10.700 2.660 10.775 3.525 ;
        RECT  4.120 2.725 10.700 3.525 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 1.790 3.030 2.130 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.080 -0.400 12.540 0.400 ;
        RECT  8.740 -0.400 9.080 0.895 ;
        RECT  7.640 -0.400 8.740 0.400 ;
        RECT  7.300 -0.400 7.640 0.895 ;
        RECT  6.320 -0.400 7.300 0.400 ;
        RECT  5.980 -0.400 6.320 0.895 ;
        RECT  5.040 -0.400 5.980 0.400 ;
        RECT  4.700 -0.400 5.040 0.895 ;
        RECT  3.760 -0.400 4.700 0.400 ;
        RECT  3.420 -0.400 3.760 0.895 ;
        RECT  2.320 -0.400 3.420 0.400 ;
        RECT  1.980 -0.400 2.320 0.895 ;
        RECT  0.000 -0.400 1.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.580 4.640 12.540 5.440 ;
        RECT  11.240 4.090 11.580 5.440 ;
        RECT  10.260 4.640 11.240 5.440 ;
        RECT  9.920 4.020 10.260 5.440 ;
        RECT  8.980 4.640 9.920 5.440 ;
        RECT  8.640 4.020 8.980 5.440 ;
        RECT  7.700 4.640 8.640 5.440 ;
        RECT  7.360 4.020 7.700 5.440 ;
        RECT  6.380 4.640 7.360 5.440 ;
        RECT  6.040 4.020 6.380 5.440 ;
        RECT  5.100 4.640 6.040 5.440 ;
        RECT  4.760 4.020 5.100 5.440 ;
        RECT  3.820 4.640 4.760 5.440 ;
        RECT  3.480 4.020 3.820 5.440 ;
        RECT  2.500 4.640 3.480 5.440 ;
        RECT  2.160 3.620 2.500 5.440 ;
        RECT  1.180 4.640 2.160 5.440 ;
        RECT  1.125 4.465 1.180 5.440 ;
        RECT  0.895 4.410 1.125 5.440 ;
        RECT  0.840 4.465 0.895 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 2.155 10.360 2.495 ;
        RECT  3.440 1.150 3.780 3.100 ;
        RECT  1.260 1.150 3.440 1.490 ;
        RECT  1.520 2.760 3.440 3.100 ;
    END
END CLKBUFX16

MACRO CLKBUFX12
    CLASS CORE ;
    FOREIGN CLKBUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.480 1.200 9.685 3.280 ;
        RECT  8.135 1.180 9.480 3.350 ;
        RECT  3.460 1.180 8.135 1.860 ;
        RECT  8.060 2.660 8.135 3.350 ;
        RECT  3.380 2.670 8.060 3.350 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.990 2.580 2.330 ;
        RECT  1.535 1.845 1.765 2.330 ;
        RECT  0.600 1.990 1.535 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.000 -0.400 10.560 0.400 ;
        RECT  6.660 -0.400 7.000 0.950 ;
        RECT  5.720 -0.400 6.660 0.400 ;
        RECT  5.380 -0.400 5.720 0.950 ;
        RECT  4.440 -0.400 5.380 0.400 ;
        RECT  4.100 -0.400 4.440 0.950 ;
        RECT  3.160 -0.400 4.100 0.400 ;
        RECT  2.820 -0.400 3.160 0.950 ;
        RECT  1.880 -0.400 2.820 0.400 ;
        RECT  1.540 -0.400 1.880 0.950 ;
        RECT  0.000 -0.400 1.540 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.520 4.640 10.560 5.440 ;
        RECT  9.465 4.465 9.520 5.440 ;
        RECT  9.235 4.410 9.465 5.440 ;
        RECT  9.180 4.465 9.235 5.440 ;
        RECT  8.200 4.640 9.180 5.440 ;
        RECT  7.860 3.675 8.200 5.440 ;
        RECT  6.920 4.640 7.860 5.440 ;
        RECT  6.580 3.675 6.920 5.440 ;
        RECT  5.640 4.640 6.580 5.440 ;
        RECT  5.300 3.675 5.640 5.440 ;
        RECT  4.360 4.640 5.300 5.440 ;
        RECT  4.020 3.675 4.360 5.440 ;
        RECT  3.080 4.640 4.020 5.440 ;
        RECT  2.740 3.725 3.080 5.440 ;
        RECT  1.800 4.640 2.740 5.440 ;
        RECT  1.460 3.705 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.705 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.150 2.090 7.800 2.430 ;
        RECT  2.810 1.340 3.150 3.100 ;
        RECT  2.180 1.340 2.810 1.680 ;
        RECT  0.820 2.760 2.810 3.100 ;
    END
END CLKBUFX12

MACRO BUFXL
    CLASS CORE ;
    FOREIGN BUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 1.150 2.425 3.050 ;
        RECT  1.880 1.150 2.195 1.380 ;
        RECT  2.120 2.635 2.195 3.050 ;
        RECT  1.840 2.820 2.120 3.050 ;
        RECT  1.540 1.040 1.880 1.380 ;
        RECT  1.500 2.820 1.840 3.160 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.810 2.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 2.640 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.270 2.060 1.520 2.400 ;
        RECT  1.040 1.220 1.270 2.990 ;
        RECT  0.520 1.220 1.040 1.450 ;
        RECT  0.520 2.760 1.040 2.990 ;
        RECT  0.180 1.110 0.520 1.450 ;
        RECT  0.180 2.760 0.520 3.100 ;
    END
END BUFXL

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.530 1.820 5.065 3.220 ;
        RECT  4.200 1.820 4.530 3.250 ;
        RECT  3.515 1.290 4.200 3.250 ;
        RECT  3.440 1.290 3.515 1.850 ;
        RECT  3.440 2.630 3.515 3.250 ;
        RECT  2.260 1.290 3.440 1.770 ;
        RECT  2.180 2.770 3.440 3.250 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 1.990 1.380 2.330 ;
        RECT  0.875 1.845 1.105 2.330 ;
        RECT  0.570 1.990 0.875 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.520 -0.400 5.940 0.400 ;
        RECT  4.180 -0.400 4.520 0.950 ;
        RECT  3.240 -0.400 4.180 0.400 ;
        RECT  2.900 -0.400 3.240 0.950 ;
        RECT  1.960 -0.400 2.900 0.400 ;
        RECT  1.620 -0.400 1.960 0.895 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 4.640 5.940 5.440 ;
        RECT  4.100 3.620 4.440 5.440 ;
        RECT  3.160 4.640 4.100 5.440 ;
        RECT  2.820 3.620 3.160 5.440 ;
        RECT  1.880 4.640 2.820 5.440 ;
        RECT  1.540 3.705 1.880 5.440 ;
        RECT  0.600 4.640 1.540 5.440 ;
        RECT  0.260 3.705 0.600 5.440 ;
        RECT  0.000 4.640 0.260 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.950 2.180 3.210 2.520 ;
        RECT  1.610 1.150 1.950 3.100 ;
        RECT  0.900 1.150 1.610 1.490 ;
        RECT  0.900 2.760 1.610 3.100 ;
    END
END BUFX8

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 1.260 2.500 3.080 ;
        RECT  2.120 1.260 2.200 3.220 ;
        RECT  2.040 1.260 2.120 1.730 ;
        RECT  2.040 2.740 2.120 3.220 ;
        RECT  1.700 0.920 2.040 1.730 ;
        RECT  1.700 2.740 2.040 4.020 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.800 2.395 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 -0.400 3.300 0.400 ;
        RECT  2.460 -0.400 2.800 0.575 ;
        RECT  1.280 -0.400 2.460 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 4.640 3.300 5.440 ;
        RECT  2.460 3.940 2.800 5.440 ;
        RECT  1.280 4.640 2.460 5.440 ;
        RECT  0.940 3.940 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.380 2.005 1.890 2.455 ;
        RECT  1.040 1.250 1.380 3.080 ;
        RECT  0.520 1.250 1.040 1.590 ;
        RECT  0.520 2.740 1.040 3.080 ;
        RECT  0.180 0.780 0.520 1.590 ;
        RECT  0.180 2.740 0.520 4.020 ;
    END
END BUFX4

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.205 1.880 1.545 ;
        RECT  1.770 1.820 1.840 3.160 ;
        RECT  1.540 1.205 1.770 3.160 ;
        RECT  1.500 1.820 1.540 3.160 ;
        RECT  1.460 1.820 1.500 2.660 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.555 2.360 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 -0.400 2.640 0.400 ;
        RECT  2.100 -0.400 2.440 0.575 ;
        RECT  0.000 -0.400 2.100 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 4.640 2.640 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.115 1.975 1.225 2.315 ;
        RECT  0.885 1.135 1.115 3.155 ;
        RECT  0.520 1.135 0.885 1.365 ;
        RECT  0.520 2.925 0.885 3.155 ;
        RECT  0.180 1.025 0.520 1.365 ;
        RECT  0.180 2.925 0.520 3.265 ;
    END
END BUFX3

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 1.845 2.425 2.075 ;
        RECT  2.120 1.500 2.350 2.980 ;
        RECT  1.980 1.500 2.120 1.730 ;
        RECT  1.940 2.750 2.120 2.980 ;
        RECT  1.640 1.390 1.980 1.730 ;
        RECT  1.600 2.750 1.940 3.090 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.890 2.260 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 -0.400 2.640 0.400 ;
        RECT  0.880 -0.400 1.220 0.575 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 2.640 5.440 ;
        RECT  1.125 4.465 1.180 5.440 ;
        RECT  0.895 4.410 1.125 5.440 ;
        RECT  0.840 4.465 0.895 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.370 2.060 1.620 2.400 ;
        RECT  1.140 1.265 1.370 2.990 ;
        RECT  0.620 1.265 1.140 1.495 ;
        RECT  0.620 2.760 1.140 2.990 ;
        RECT  0.280 1.155 0.620 1.495 ;
        RECT  0.280 2.760 0.620 3.100 ;
    END
END BUFX2

MACRO BUFX20
    CLASS CORE ;
    FOREIGN BUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.795 1.125 10.345 3.840 ;
        RECT  3.420 1.125 8.795 1.925 ;
        RECT  8.720 2.660 8.795 3.525 ;
        RECT  3.380 2.725 8.720 3.525 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.990 2.500 2.330 ;
        RECT  1.535 1.845 1.765 2.330 ;
        RECT  0.750 1.990 1.535 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.560 -0.400 10.560 0.400 ;
        RECT  9.220 -0.400 9.560 0.575 ;
        RECT  8.240 -0.400 9.220 0.400 ;
        RECT  7.900 -0.400 8.240 0.895 ;
        RECT  6.960 -0.400 7.900 0.400 ;
        RECT  6.620 -0.400 6.960 0.895 ;
        RECT  5.680 -0.400 6.620 0.400 ;
        RECT  5.340 -0.400 5.680 0.895 ;
        RECT  4.400 -0.400 5.340 0.400 ;
        RECT  4.060 -0.400 4.400 0.895 ;
        RECT  3.120 -0.400 4.060 0.400 ;
        RECT  2.780 -0.400 3.120 0.965 ;
        RECT  1.800 -0.400 2.780 0.400 ;
        RECT  1.460 -0.400 1.800 1.045 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 1.045 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.520 4.640 10.560 5.440 ;
        RECT  9.465 4.465 9.520 5.440 ;
        RECT  9.235 4.410 9.465 5.440 ;
        RECT  9.180 4.465 9.235 5.440 ;
        RECT  8.200 4.640 9.180 5.440 ;
        RECT  7.860 4.090 8.200 5.440 ;
        RECT  6.920 4.640 7.860 5.440 ;
        RECT  6.580 4.090 6.920 5.440 ;
        RECT  5.640 4.640 6.580 5.440 ;
        RECT  5.300 4.020 5.640 5.440 ;
        RECT  4.360 4.640 5.300 5.440 ;
        RECT  4.020 4.020 4.360 5.440 ;
        RECT  3.080 4.640 4.020 5.440 ;
        RECT  2.740 3.605 3.080 5.440 ;
        RECT  1.800 4.640 2.740 5.440 ;
        RECT  1.460 3.605 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.605 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.145 2.155 8.260 2.495 ;
        RECT  2.805 1.345 3.145 3.180 ;
        RECT  2.100 1.345 2.805 1.685 ;
        RECT  0.820 2.840 2.805 3.180 ;
        RECT  1.160 1.345 2.100 1.575 ;
        RECT  0.820 1.345 1.160 1.685 ;
    END
END BUFX20

MACRO BUFX1
    CLASS CORE ;
    FOREIGN BUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 1.150 2.425 3.050 ;
        RECT  1.880 1.150 2.195 1.380 ;
        RECT  2.120 2.635 2.195 3.050 ;
        RECT  1.840 2.820 2.120 3.050 ;
        RECT  1.540 1.040 1.880 1.380 ;
        RECT  1.500 2.820 1.840 3.160 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.810 2.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 -0.400 2.640 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 2.640 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.270 2.060 1.520 2.400 ;
        RECT  1.040 1.220 1.270 2.990 ;
        RECT  0.520 1.220 1.040 1.450 ;
        RECT  0.520 2.760 1.040 2.990 ;
        RECT  0.180 1.110 0.520 1.450 ;
        RECT  0.180 2.760 0.520 3.100 ;
    END
END BUFX1

MACRO BUFX16
    CLASS CORE ;
    FOREIGN BUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.125 8.365 3.840 ;
        RECT  2.780 1.125 6.815 1.925 ;
        RECT  6.740 2.625 6.815 3.525 ;
        RECT  3.420 2.725 6.740 3.525 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 2.190 2.040 2.530 ;
        RECT  1.535 2.190 1.765 2.635 ;
        RECT  0.580 2.190 1.535 2.530 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.720 -0.400 8.580 0.400 ;
        RECT  7.380 -0.400 7.720 0.575 ;
        RECT  6.360 -0.400 7.380 0.400 ;
        RECT  6.020 -0.400 6.360 0.895 ;
        RECT  5.040 -0.400 6.020 0.400 ;
        RECT  4.700 -0.400 5.040 0.895 ;
        RECT  3.760 -0.400 4.700 0.400 ;
        RECT  3.420 -0.400 3.760 0.895 ;
        RECT  2.440 -0.400 3.420 0.400 ;
        RECT  2.100 -0.400 2.440 0.970 ;
        RECT  1.160 -0.400 2.100 0.400 ;
        RECT  0.820 -0.400 1.160 0.965 ;
        RECT  0.000 -0.400 0.820 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.400 4.640 8.580 5.440 ;
        RECT  8.060 4.465 8.400 5.440 ;
        RECT  7.040 4.640 8.060 5.440 ;
        RECT  6.700 4.465 7.040 5.440 ;
        RECT  5.680 4.640 6.700 5.440 ;
        RECT  5.340 4.020 5.680 5.440 ;
        RECT  4.400 4.640 5.340 5.440 ;
        RECT  4.060 4.020 4.400 5.440 ;
        RECT  3.120 4.640 4.060 5.440 ;
        RECT  2.780 4.020 3.120 5.440 ;
        RECT  1.800 4.640 2.780 5.440 ;
        RECT  1.460 3.395 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.395 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.505 2.155 6.510 2.495 ;
        RECT  2.275 1.405 2.505 3.120 ;
        RECT  0.180 1.405 2.275 1.745 ;
        RECT  2.100 2.760 2.275 3.120 ;
        RECT  1.160 2.890 2.100 3.120 ;
        RECT  0.820 2.760 1.160 3.120 ;
    END
END BUFX16

MACRO BUFX12
    CLASS CORE ;
    FOREIGN BUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.260 6.385 3.220 ;
        RECT  4.760 1.350 4.835 1.850 ;
        RECT  4.760 2.630 4.835 3.180 ;
        RECT  2.820 1.350 4.760 1.690 ;
        RECT  2.740 2.840 4.760 3.180 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 1.990 2.030 2.330 ;
        RECT  0.875 1.845 1.105 2.330 ;
        RECT  0.710 1.990 0.875 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.360 -0.400 6.600 0.400 ;
        RECT  6.020 -0.400 6.360 0.950 ;
        RECT  5.080 -0.400 6.020 0.400 ;
        RECT  4.740 -0.400 5.080 0.950 ;
        RECT  3.800 -0.400 4.740 0.400 ;
        RECT  3.460 -0.400 3.800 0.965 ;
        RECT  2.520 -0.400 3.460 0.400 ;
        RECT  2.180 -0.400 2.520 0.965 ;
        RECT  1.200 -0.400 2.180 0.400 ;
        RECT  0.860 -0.400 1.200 0.575 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 4.640 6.600 5.440 ;
        RECT  6.080 4.020 6.420 5.440 ;
        RECT  5.050 4.640 6.080 5.440 ;
        RECT  4.710 4.020 5.050 5.440 ;
        RECT  3.720 4.640 4.710 5.440 ;
        RECT  3.380 4.020 3.720 5.440 ;
        RECT  2.440 4.640 3.380 5.440 ;
        RECT  2.100 3.705 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 3.705 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.510 2.180 4.375 2.520 ;
        RECT  2.280 1.450 2.510 2.990 ;
        RECT  1.880 1.450 2.280 1.680 ;
        RECT  1.800 2.760 2.280 2.990 ;
        RECT  1.540 1.340 1.880 1.680 ;
        RECT  1.460 2.760 1.800 3.100 ;
        RECT  0.520 1.340 1.540 1.570 ;
        RECT  0.520 2.760 1.460 2.990 ;
        RECT  0.290 1.340 0.520 1.635 ;
        RECT  0.180 2.760 0.520 3.100 ;
        RECT  0.180 1.405 0.290 1.635 ;
    END
END BUFX12

MACRO AOI33XL
    CLASS CORE ;
    FOREIGN AOI33XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.240 5.065 3.450 ;
        RECT  2.110 1.240 4.835 1.470 ;
        RECT  4.560 3.220 4.835 3.450 ;
        RECT  4.220 3.220 4.560 3.560 ;
        RECT  3.120 3.220 4.220 3.450 ;
        RECT  2.780 3.220 3.120 3.560 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.685 0.630 2.195 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 2.685 1.410 3.025 ;
        RECT  0.755 2.685 1.290 3.195 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.580 1.700 2.090 2.125 ;
        RECT  1.535 1.845 1.580 2.075 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.050 1.715 4.480 2.215 ;
        RECT  3.980 1.715 4.050 2.120 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 2.265 3.745 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.170 2.405 2.710 2.940 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 -0.400 5.280 0.400 ;
        RECT  3.990 -0.400 4.330 0.575 ;
        RECT  0.520 -0.400 3.990 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 4.640 5.280 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.520 4.640 1.300 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.460 3.695 3.840 4.025 ;
        RECT  2.400 3.795 3.460 4.025 ;
        RECT  2.115 3.640 2.400 4.025 ;
        RECT  0.740 3.640 2.115 3.980 ;
    END
END AOI33XL

MACRO AOI33X4
    CLASS CORE ;
    FOREIGN AOI33X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI33XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.970 1.820 7.120 3.220 ;
        RECT  6.740 1.430 6.970 3.220 ;
        RECT  6.405 1.430 6.740 1.660 ;
        RECT  6.065 2.820 6.740 3.160 ;
        RECT  6.065 1.320 6.405 1.660 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.650 0.615 2.100 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.355 1.425 2.905 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.750 2.160 2.100 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.055 2.105 4.480 2.660 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 1.820 3.820 2.150 ;
        RECT  2.970 1.920 2.975 2.150 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 2.405 3.160 2.880 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 -0.400 7.260 0.400 ;
        RECT  6.705 -0.400 7.045 0.960 ;
        RECT  5.725 -0.400 6.705 0.400 ;
        RECT  5.385 -0.400 5.725 0.900 ;
        RECT  4.280 -0.400 5.385 0.400 ;
        RECT  3.940 -0.400 4.280 0.575 ;
        RECT  0.520 -0.400 3.940 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 4.640 7.260 5.440 ;
        RECT  6.705 3.680 7.045 5.440 ;
        RECT  5.765 4.640 6.705 5.440 ;
        RECT  5.425 3.870 5.765 5.440 ;
        RECT  1.645 4.640 5.425 5.440 ;
        RECT  1.305 4.465 1.645 5.440 ;
        RECT  0.525 4.640 1.305 5.440 ;
        RECT  0.185 4.465 0.525 5.440 ;
        RECT  0.000 4.640 0.185 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.430 2.085 6.440 2.315 ;
        RECT  5.200 1.180 5.430 3.585 ;
        RECT  5.010 1.180 5.200 1.410 ;
        RECT  5.110 3.355 5.200 3.585 ;
        RECT  4.880 3.355 5.110 4.045 ;
        RECT  4.780 0.665 5.010 1.410 ;
        RECT  4.725 1.645 4.955 3.120 ;
        RECT  4.665 3.815 4.880 4.045 ;
        RECT  4.665 0.665 4.780 0.895 ;
        RECT  4.285 1.645 4.725 1.875 ;
        RECT  4.405 2.890 4.725 3.120 ;
        RECT  4.175 2.890 4.405 3.370 ;
        RECT  4.055 1.160 4.285 1.875 ;
        RECT  3.070 3.140 4.175 3.370 ;
        RECT  2.345 1.160 4.055 1.390 ;
        RECT  3.545 3.925 3.895 4.405 ;
        RECT  2.350 3.925 3.545 4.155 ;
        RECT  2.840 3.140 3.070 3.525 ;
        RECT  2.120 3.265 2.350 4.155 ;
        RECT  2.115 1.025 2.345 1.390 ;
        RECT  0.800 3.265 2.120 3.605 ;
    END
END AOI33X4

MACRO AOI33X2
    CLASS CORE ;
    FOREIGN AOI33X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI33XL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.135 0.805 8.365 3.305 ;
        RECT  8.060 0.805 8.135 1.285 ;
        RECT  4.745 3.075 8.135 3.305 ;
        RECT  3.530 0.805 8.060 1.035 ;
        RECT  3.300 0.805 3.530 1.480 ;
        RECT  2.020 1.250 3.300 1.480 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 2.850 3.995 3.190 ;
        RECT  0.700 2.960 3.615 3.190 ;
        RECT  0.470 2.405 0.700 3.190 ;
        RECT  0.215 2.405 0.470 2.635 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.500 3.275 2.730 ;
        RECT  2.855 1.845 3.085 2.730 ;
        RECT  1.095 2.500 2.855 2.730 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 1.845 2.155 2.270 ;
        RECT  1.535 1.845 1.780 2.075 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.600 1.265 7.830 2.020 ;
        RECT  4.470 1.265 7.600 1.495 ;
        RECT  4.240 1.265 4.470 2.325 ;
        RECT  4.175 1.845 4.240 2.075 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.770 1.725 7.000 2.410 ;
        RECT  5.270 1.725 6.770 1.955 ;
        RECT  5.040 1.725 5.270 2.690 ;
        RECT  4.835 2.405 5.040 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.750 2.205 6.460 2.660 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.005 -0.400 8.580 0.400 ;
        RECT  7.665 -0.400 8.005 0.575 ;
        RECT  4.245 -0.400 7.665 0.400 ;
        RECT  3.905 -0.400 4.245 0.575 ;
        RECT  0.520 -0.400 3.905 0.400 ;
        RECT  0.180 -0.400 0.520 1.755 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 4.640 8.580 5.440 ;
        RECT  3.380 4.070 3.720 5.440 ;
        RECT  2.440 4.640 3.380 5.440 ;
        RECT  2.100 4.070 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 4.070 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.955 3.765 8.295 4.105 ;
        RECT  7.005 3.820 7.955 4.050 ;
        RECT  6.665 3.765 7.005 4.105 ;
        RECT  5.725 3.820 6.665 4.050 ;
        RECT  5.385 3.765 5.725 4.105 ;
        RECT  4.445 3.820 5.385 4.050 ;
        RECT  4.335 3.765 4.445 4.105 ;
        RECT  4.105 3.420 4.335 4.105 ;
        RECT  0.180 3.420 4.105 3.650 ;
    END
END AOI33X2

MACRO AOI33X1
    CLASS CORE ;
    FOREIGN AOI33X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI33XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.990 2.405 5.065 2.635 ;
        RECT  4.835 0.905 4.990 3.135 ;
        RECT  4.760 0.905 4.835 3.220 ;
        RECT  2.020 0.905 4.760 1.135 ;
        RECT  4.720 2.905 4.760 3.220 ;
        RECT  4.380 2.905 4.720 3.830 ;
        RECT  3.515 2.905 4.380 3.135 ;
        RECT  2.940 2.905 3.515 3.245 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.760 0.840 2.145 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 2.380 1.475 2.770 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.420 1.660 2.135 2.100 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.900 1.610 4.405 2.130 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 2.380 3.915 2.660 ;
        RECT  3.180 2.295 3.520 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.410 2.295 2.925 2.660 ;
        RECT  2.195 2.405 2.410 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.240 -0.400 5.280 0.400 ;
        RECT  3.900 -0.400 4.240 0.575 ;
        RECT  0.520 -0.400 3.900 0.400 ;
        RECT  0.180 -0.400 0.520 1.430 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 4.640 5.280 5.440 ;
        RECT  1.660 4.465 2.000 5.440 ;
        RECT  0.520 4.640 1.660 5.440 ;
        RECT  0.180 3.010 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.660 3.610 4.000 4.005 ;
        RECT  2.560 3.775 3.660 4.005 ;
        RECT  2.220 3.010 2.560 4.005 ;
        RECT  1.240 3.775 2.220 4.005 ;
        RECT  0.900 3.010 1.240 4.005 ;
    END
END AOI33X1

MACRO AOI32XL
    CLASS CORE ;
    FOREIGN AOI32XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 1.845 4.405 2.075 ;
        RECT  4.100 1.455 4.330 3.315 ;
        RECT  2.305 1.455 4.100 1.685 ;
        RECT  3.400 3.085 4.100 3.315 ;
        RECT  3.170 3.085 3.400 3.685 ;
        RECT  3.060 3.345 3.170 3.685 ;
        RECT  2.075 1.075 2.305 1.685 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.390 2.185 3.820 2.720 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.580 2.265 3.085 2.785 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.760 2.130 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.405 1.560 2.910 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.920 2.120 2.150 ;
        RECT  1.240 1.820 1.840 2.150 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.640 -0.400 4.620 0.400 ;
        RECT  3.300 -0.400 3.640 1.220 ;
        RECT  0.520 -0.400 3.300 0.400 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 4.640 4.620 5.440 ;
        RECT  1.620 3.765 1.960 5.440 ;
        RECT  0.520 4.640 1.620 5.440 ;
        RECT  0.180 3.555 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 3.640 4.120 4.145 ;
        RECT  2.680 3.915 3.780 4.145 ;
        RECT  2.340 3.300 2.680 4.145 ;
        RECT  1.240 3.300 2.340 3.530 ;
        RECT  0.900 3.300 1.240 3.895 ;
    END
END AOI32XL

MACRO AOI32X4
    CLASS CORE ;
    FOREIGN AOI32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI32XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 1.820 6.460 3.220 ;
        RECT  6.080 1.500 6.310 3.220 ;
        RECT  5.775 1.500 6.080 1.730 ;
        RECT  5.415 2.740 6.080 3.080 ;
        RECT  5.435 1.390 5.775 1.730 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.585 2.380 3.785 3.080 ;
        RECT  3.350 2.175 3.585 3.080 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.380 2.630 2.955 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.575 0.765 2.100 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.495 2.885 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.725 2.075 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 -0.400 6.600 0.400 ;
        RECT  6.080 -0.400 6.420 0.955 ;
        RECT  5.080 -0.400 6.080 0.400 ;
        RECT  4.850 -0.400 5.080 0.950 ;
        RECT  3.680 -0.400 4.850 0.400 ;
        RECT  3.340 -0.400 3.680 0.575 ;
        RECT  0.520 -0.400 3.340 0.400 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.395 4.640 6.600 5.440 ;
        RECT  6.055 3.705 6.395 5.440 ;
        RECT  5.110 4.640 6.055 5.440 ;
        RECT  4.770 3.705 5.110 5.440 ;
        RECT  1.780 4.640 4.770 5.440 ;
        RECT  1.440 4.465 1.780 5.440 ;
        RECT  0.535 4.640 1.440 5.440 ;
        RECT  0.150 4.465 0.535 5.440 ;
        RECT  0.000 4.640 0.150 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.040 2.060 5.845 2.400 ;
        RECT  4.810 1.270 5.040 3.165 ;
        RECT  4.550 1.270 4.810 1.500 ;
        RECT  4.385 2.935 4.810 3.165 ;
        RECT  4.520 1.860 4.575 2.200 ;
        RECT  4.320 0.665 4.550 1.500 ;
        RECT  4.235 1.855 4.520 2.200 ;
        RECT  4.045 2.880 4.385 3.220 ;
        RECT  4.075 0.665 4.320 0.895 ;
        RECT  4.055 1.855 4.235 2.145 ;
        RECT  3.825 1.125 4.055 2.145 ;
        RECT  3.735 3.585 3.845 3.925 ;
        RECT  3.120 1.125 3.825 1.355 ;
        RECT  3.505 3.585 3.735 4.330 ;
        RECT  2.405 4.100 3.505 4.330 ;
        RECT  3.120 3.385 3.125 3.725 ;
        RECT  2.890 1.125 3.120 3.725 ;
        RECT  2.360 1.125 2.890 1.355 ;
        RECT  2.785 3.385 2.890 3.725 ;
        RECT  2.175 3.385 2.405 4.330 ;
        RECT  2.020 1.015 2.360 1.355 ;
        RECT  2.065 3.385 2.175 3.725 ;
        RECT  1.080 3.440 2.065 3.670 ;
        RECT  0.740 3.385 1.080 3.725 ;
    END
END AOI32X4

MACRO AOI32X2
    CLASS CORE ;
    FOREIGN AOI32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI32XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.460 7.045 3.315 ;
        RECT  6.740 1.460 6.815 1.845 ;
        RECT  6.375 3.085 6.815 3.315 ;
        RECT  6.270 1.460 6.740 1.690 ;
        RECT  6.035 3.030 6.375 3.370 ;
        RECT  6.040 1.180 6.270 1.690 ;
        RECT  3.245 1.180 6.040 1.410 ;
        RECT  5.095 3.075 6.035 3.305 ;
        RECT  4.755 3.020 5.095 3.360 ;
        RECT  3.015 0.795 3.245 1.410 ;
        RECT  2.020 0.795 3.015 1.025 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.505 2.545 6.325 2.775 ;
        RECT  4.275 1.845 4.505 2.775 ;
        RECT  4.175 1.845 4.275 2.130 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.320 1.820 5.800 2.130 ;
        RECT  4.980 1.820 5.320 2.310 ;
        RECT  4.975 1.820 4.980 2.130 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.605 2.390 3.835 2.905 ;
        RECT  3.440 2.630 3.605 2.905 ;
        RECT  0.645 2.675 3.440 2.905 ;
        RECT  0.415 2.405 0.645 2.905 ;
        RECT  0.215 2.405 0.415 2.635 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.845 3.165 2.425 ;
        RECT  1.095 2.195 2.780 2.425 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 1.735 2.120 1.965 ;
        RECT  1.780 1.285 2.010 1.965 ;
        RECT  1.535 1.285 1.780 1.515 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.840 -0.400 7.260 0.400 ;
        RECT  6.500 -0.400 6.840 1.220 ;
        RECT  4.240 -0.400 6.500 0.400 ;
        RECT  3.900 -0.400 4.240 0.575 ;
        RECT  0.465 -0.400 3.900 0.400 ;
        RECT  0.235 -0.400 0.465 1.430 ;
        RECT  0.000 -0.400 0.235 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.725 4.640 7.260 5.440 ;
        RECT  3.385 4.090 3.725 5.440 ;
        RECT  2.445 4.640 3.385 5.440 ;
        RECT  2.105 4.090 2.445 5.440 ;
        RECT  1.160 4.640 2.105 5.440 ;
        RECT  0.820 4.090 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.675 3.765 7.015 4.105 ;
        RECT  5.735 3.820 6.675 4.050 ;
        RECT  5.395 3.765 5.735 4.105 ;
        RECT  4.455 3.820 5.395 4.050 ;
        RECT  4.345 3.765 4.455 4.105 ;
        RECT  4.115 3.410 4.345 4.105 ;
        RECT  3.085 3.410 4.115 3.640 ;
        RECT  2.745 3.355 3.085 3.695 ;
        RECT  1.805 3.400 2.745 3.630 ;
        RECT  1.465 3.345 1.805 3.685 ;
        RECT  0.520 3.400 1.465 3.630 ;
        RECT  0.180 3.345 0.520 3.685 ;
    END
END AOI32X2

MACRO AOI32X1
    CLASS CORE ;
    FOREIGN AOI32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI32XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 0.935 4.405 3.445 ;
        RECT  4.100 0.935 4.175 1.285 ;
        RECT  3.060 3.215 4.175 3.445 ;
        RECT  2.020 0.935 4.100 1.165 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.115 1.600 3.745 2.075 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.530 2.350 3.160 2.690 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.800 2.100 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.400 1.480 2.855 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.610 2.120 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.710 -0.400 4.620 0.400 ;
        RECT  3.370 -0.400 3.710 0.575 ;
        RECT  0.465 -0.400 3.370 0.400 ;
        RECT  0.235 -0.400 0.465 1.430 ;
        RECT  0.000 -0.400 0.235 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 4.640 4.620 5.440 ;
        RECT  1.620 3.820 1.960 5.440 ;
        RECT  0.520 4.640 1.620 5.440 ;
        RECT  0.180 3.295 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.625 3.815 4.120 4.045 ;
        RECT  2.395 3.360 2.625 4.045 ;
        RECT  0.900 3.360 2.395 3.590 ;
    END
END AOI32X1

MACRO AOI31XL
    CLASS CORE ;
    FOREIGN AOI31XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 1.175 3.085 1.515 ;
        RECT  2.835 1.175 3.065 3.320 ;
        RECT  2.020 1.175 2.835 1.405 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 2.375 2.585 2.755 ;
        RECT  1.960 2.380 2.355 2.755 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.600 0.520 2.185 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.485 2.730 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.640 2.280 2.100 ;
        RECT  1.535 1.845 1.540 2.075 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 -0.400 3.300 0.400 ;
        RECT  2.725 -0.400 3.065 0.575 ;
        RECT  0.520 -0.400 2.725 0.400 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 4.640 3.300 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.545 4.640 1.500 5.440 ;
        RECT  0.175 4.465 0.545 5.440 ;
        RECT  0.000 4.640 0.175 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.740 3.190 2.400 3.530 ;
    END
END AOI31XL

MACRO AOI31X4
    CLASS CORE ;
    FOREIGN AOI31X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI31XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.820 5.800 3.220 ;
        RECT  5.420 1.415 5.740 3.220 ;
        RECT  4.685 1.415 5.420 1.645 ;
        RECT  4.690 2.800 5.420 3.030 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 1.800 3.160 2.370 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.525 0.520 2.100 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 2.380 1.265 3.050 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.415 1.720 1.935 2.130 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.670 -0.400 5.940 0.400 ;
        RECT  5.330 -0.400 5.670 0.960 ;
        RECT  4.385 -0.400 5.330 0.400 ;
        RECT  4.045 -0.400 4.385 0.960 ;
        RECT  2.960 -0.400 4.045 0.400 ;
        RECT  2.620 -0.400 2.960 0.575 ;
        RECT  0.520 -0.400 2.620 0.400 ;
        RECT  0.180 -0.400 0.520 1.290 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 4.640 5.940 5.440 ;
        RECT  5.385 3.735 5.615 5.440 ;
        RECT  4.385 4.640 5.385 5.440 ;
        RECT  4.045 3.760 4.385 5.440 ;
        RECT  1.640 4.640 4.045 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.520 4.640 1.300 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.090 2.035 5.185 2.400 ;
        RECT  3.860 1.315 4.090 3.435 ;
        RECT  3.605 1.315 3.860 1.545 ;
        RECT  3.680 3.205 3.860 3.435 ;
        RECT  3.450 3.205 3.680 4.375 ;
        RECT  3.390 1.860 3.620 2.930 ;
        RECT  3.375 0.640 3.605 1.545 ;
        RECT  3.325 4.145 3.450 4.375 ;
        RECT  3.065 2.700 3.390 2.930 ;
        RECT  2.835 2.700 3.065 3.640 ;
        RECT  2.395 2.700 2.835 2.930 ;
        RECT  0.740 3.525 2.400 3.755 ;
        RECT  2.165 1.115 2.395 2.930 ;
        RECT  2.075 1.115 2.165 1.485 ;
    END
END AOI31X4

MACRO AOI31X2
    CLASS CORE ;
    FOREIGN AOI31X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI31XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.795 2.635 5.025 3.360 ;
        RECT  4.760 2.635 4.795 2.965 ;
        RECT  4.405 2.635 4.760 2.865 ;
        RECT  4.175 1.125 4.405 2.865 ;
        RECT  1.790 1.125 4.175 1.355 ;
        RECT  1.560 0.665 1.790 1.355 ;
        RECT  0.180 0.665 1.560 0.895 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.635 1.820 5.180 2.340 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.735 2.280 1.965 ;
        RECT  0.875 1.285 1.180 1.965 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.160 2.215 3.275 2.445 ;
        RECT  2.780 1.845 3.160 2.445 ;
        RECT  1.220 2.215 2.780 2.445 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 2.060 3.905 2.905 ;
        RECT  0.520 2.675 3.675 2.905 ;
        RECT  0.140 2.310 0.520 2.905 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.960 -0.400 5.940 0.400 ;
        RECT  4.940 -0.400 4.960 0.575 ;
        RECT  4.710 -0.400 4.940 1.340 ;
        RECT  4.620 -0.400 4.710 0.575 ;
        RECT  2.360 -0.400 4.620 0.400 ;
        RECT  2.020 -0.400 2.360 0.895 ;
        RECT  0.000 -0.400 2.020 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 4.640 5.940 5.440 ;
        RECT  3.380 3.765 3.720 5.440 ;
        RECT  2.440 4.640 3.380 5.440 ;
        RECT  2.100 3.765 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 3.765 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.190 3.820 5.720 4.050 ;
        RECT  3.960 3.135 4.190 4.050 ;
        RECT  0.180 3.135 3.960 3.365 ;
    END
END AOI31X2

MACRO AOI31X1
    CLASS CORE ;
    FOREIGN AOI31X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI31XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.025 0.845 3.085 3.175 ;
        RECT  2.855 0.845 3.025 4.025 ;
        RECT  2.780 0.845 2.855 1.540 ;
        RECT  2.795 2.945 2.855 4.025 ;
        RECT  2.020 0.845 2.780 1.075 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.620 2.105 2.625 2.450 ;
        RECT  2.230 2.105 2.620 2.660 ;
        RECT  2.120 2.380 2.230 2.660 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.765 0.520 2.400 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.345 1.295 2.805 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.670 1.940 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 -0.400 3.300 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  0.520 -0.400 2.780 0.400 ;
        RECT  0.180 -0.400 0.520 0.895 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 4.640 3.300 5.440 ;
        RECT  1.460 3.780 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.785 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.820 3.040 2.440 3.270 ;
    END
END AOI31X1

MACRO AOI2BB2XL
    CLASS CORE ;
    FOREIGN AOI2BB2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.430 4.205 3.555 ;
        RECT  3.745 2.430 3.975 2.660 ;
        RECT  3.515 1.275 3.745 2.660 ;
        RECT  3.090 1.275 3.515 1.505 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.135 2.380 2.500 2.965 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 1.885 3.160 2.660 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.590 0.755 2.100 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.495 1.180 3.220 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 -0.400 4.620 0.400 ;
        RECT  3.760 -0.400 4.100 0.575 ;
        RECT  2.120 -0.400 3.760 0.400 ;
        RECT  1.780 -0.400 2.120 0.575 ;
        RECT  0.520 -0.400 1.780 0.400 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 4.640 4.620 5.440 ;
        RECT  2.440 4.465 2.780 5.440 ;
        RECT  0.520 4.640 2.440 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.975 0.810 4.205 2.095 ;
        RECT  1.640 0.810 3.975 1.040 ;
        RECT  3.200 3.635 3.540 3.975 ;
        RECT  2.165 3.690 3.200 3.920 ;
        RECT  1.935 3.215 2.165 3.920 ;
        RECT  1.410 0.810 1.640 4.280 ;
        RECT  0.980 0.990 1.410 1.220 ;
        RECT  1.395 3.920 1.410 4.280 ;
    END
END AOI2BB2XL

MACRO AOI2BB2X4
    CLASS CORE ;
    FOREIGN AOI2BB2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB2XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 0.700 8.440 2.100 ;
        RECT  3.535 1.130 8.060 1.360 ;
        RECT  3.520 4.110 4.740 4.340 ;
        RECT  3.520 0.930 3.535 1.360 ;
        RECT  3.290 0.930 3.520 4.340 ;
        RECT  3.120 4.110 3.290 4.340 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 2.465 8.740 2.695 ;
        RECT  7.435 1.840 7.665 2.695 ;
        RECT  5.065 1.840 7.435 2.070 ;
        RECT  4.495 1.840 5.065 2.075 ;
        RECT  4.265 1.840 4.495 2.325 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.955 2.380 6.460 2.805 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 2.965 2.425 3.195 ;
        RECT  1.915 1.930 2.145 4.165 ;
        RECT  0.520 3.935 1.915 4.165 ;
        RECT  0.475 3.755 0.520 4.165 ;
        RECT  0.245 2.360 0.475 4.165 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 1.715 1.220 2.210 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.095 -0.400 9.900 0.400 ;
        RECT  6.755 -0.400 7.095 0.895 ;
        RECT  4.310 -0.400 6.755 0.400 ;
        RECT  3.970 -0.400 4.310 0.895 ;
        RECT  2.485 -0.400 3.970 0.400 ;
        RECT  2.145 -0.400 2.485 0.575 ;
        RECT  0.915 -0.400 2.145 0.400 ;
        RECT  0.575 -0.400 0.915 0.895 ;
        RECT  0.000 -0.400 0.575 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.580 4.640 9.900 5.440 ;
        RECT  8.240 4.055 8.580 5.440 ;
        RECT  7.300 4.640 8.240 5.440 ;
        RECT  6.960 4.055 7.300 5.440 ;
        RECT  6.020 4.640 6.960 5.440 ;
        RECT  5.680 4.055 6.020 5.440 ;
        RECT  2.760 4.640 5.680 5.440 ;
        RECT  2.420 4.465 2.760 5.440 ;
        RECT  0.520 4.640 2.420 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.760 3.095 9.220 3.325 ;
        RECT  2.825 1.135 3.055 2.260 ;
        RECT  1.680 1.135 2.825 1.365 ;
        RECT  1.450 1.135 1.680 3.295 ;
        RECT  1.365 1.135 1.450 1.365 ;
        RECT  1.355 2.930 1.450 3.295 ;
    END
END AOI2BB2X4

MACRO AOI2BB2X2
    CLASS CORE ;
    FOREIGN AOI2BB2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB2XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.600 1.285 5.725 1.515 ;
        RECT  5.370 0.805 5.600 4.105 ;
        RECT  2.870 0.805 5.370 1.035 ;
        RECT  4.840 3.875 5.370 4.105 ;
        RECT  4.465 3.875 4.840 4.370 ;
        RECT  4.405 4.060 4.465 4.370 ;
        RECT  4.060 4.140 4.405 4.370 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 2.280 4.460 3.095 ;
        RECT  1.900 2.865 4.100 3.095 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 1.590 5.090 2.090 ;
        RECT  2.495 1.590 4.805 1.820 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 1.630 1.840 2.100 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.870 0.520 2.660 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 -0.400 5.940 0.400 ;
        RECT  3.640 -0.400 3.980 0.575 ;
        RECT  1.915 -0.400 3.640 0.400 ;
        RECT  1.575 -0.400 1.915 1.275 ;
        RECT  0.520 -0.400 1.575 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 4.640 5.940 5.440 ;
        RECT  5.380 4.465 5.720 5.440 ;
        RECT  3.120 4.640 5.380 5.440 ;
        RECT  2.780 4.085 3.120 5.440 ;
        RECT  1.840 4.640 2.780 5.440 ;
        RECT  1.500 4.085 1.840 5.440 ;
        RECT  0.000 4.640 1.500 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.140 3.395 5.040 3.625 ;
        RECT  1.025 2.400 3.680 2.630 ;
        RECT  0.795 1.210 1.025 3.310 ;
        RECT  0.180 3.080 0.795 3.310 ;
    END
END AOI2BB2X2

MACRO AOI2BB2X1
    CLASS CORE ;
    FOREIGN AOI2BB2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.900 1.115 4.130 4.405 ;
        RECT  2.700 1.115 3.900 1.345 ;
        RECT  3.515 2.380 3.900 2.660 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 2.775 2.500 3.220 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 2.250 3.085 2.635 ;
        RECT  2.620 2.250 2.855 2.480 ;
        RECT  2.390 2.105 2.620 2.480 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.190 1.820 0.475 2.605 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 2.250 1.235 2.735 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.800 -0.400 4.620 0.400 ;
        RECT  3.460 -0.400 3.800 0.575 ;
        RECT  1.720 -0.400 3.460 0.400 ;
        RECT  1.380 -0.400 1.720 0.575 ;
        RECT  0.520 -0.400 1.380 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.900 4.640 4.620 5.440 ;
        RECT  2.560 4.090 2.900 5.440 ;
        RECT  0.520 4.640 2.560 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.290 3.450 3.540 3.680 ;
        RECT  3.235 1.575 3.465 1.990 ;
        RECT  1.700 1.575 3.235 1.805 ;
        RECT  2.060 3.450 2.290 4.375 ;
        RECT  1.840 4.145 2.060 4.375 ;
        RECT  1.470 1.575 1.700 3.420 ;
        RECT  1.065 1.575 1.470 1.805 ;
        RECT  1.355 3.050 1.470 3.420 ;
        RECT  0.835 1.315 1.065 1.805 ;
    END
END AOI2BB2X1

MACRO AOI2BB1XL
    CLASS CORE ;
    FOREIGN AOI2BB1XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.905 3.525 3.085 3.755 ;
        RECT  2.675 1.620 2.905 3.810 ;
        RECT  2.105 1.620 2.675 1.850 ;
        RECT  1.875 1.460 2.105 1.850 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.670 1.950 3.220 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.260 1.105 2.635 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.175 2.895 0.730 3.315 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 -0.400 3.300 0.400 ;
        RECT  0.930 -0.400 1.270 0.575 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 4.640 3.300 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.000 4.640 1.300 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.180 2.085 2.410 3.785 ;
        RECT  1.640 2.085 2.180 2.315 ;
        RECT  0.180 3.555 2.180 3.785 ;
        RECT  1.410 1.315 1.640 2.315 ;
        RECT  0.450 1.315 1.410 1.545 ;
    END
END AOI2BB1XL

MACRO AOI2BB1X4
    CLASS CORE ;
    FOREIGN AOI2BB1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB1XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.160 2.965 6.440 3.195 ;
        RECT  5.875 2.940 6.160 3.220 ;
        RECT  5.800 1.335 5.875 3.755 ;
        RECT  5.645 1.335 5.800 4.340 ;
        RECT  4.165 1.335 5.645 1.565 ;
        RECT  5.420 2.940 5.645 4.340 ;
        RECT  3.700 2.965 5.420 3.195 ;
        RECT  3.935 1.335 4.165 1.730 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.820 3.240 2.530 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.385 1.845 2.425 2.075 ;
        RECT  2.155 1.845 2.385 3.735 ;
        RECT  0.475 3.505 2.155 3.735 ;
        RECT  0.245 2.380 0.475 3.735 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.985 1.845 1.215 2.720 ;
        RECT  0.875 1.845 0.985 2.075 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.520 -0.400 7.260 0.400 ;
        RECT  6.180 -0.400 6.520 0.575 ;
        RECT  4.940 -0.400 6.180 0.400 ;
        RECT  4.600 -0.400 4.940 0.895 ;
        RECT  3.465 -0.400 4.600 0.400 ;
        RECT  3.125 -0.400 3.465 0.895 ;
        RECT  2.040 -0.400 3.125 0.400 ;
        RECT  1.700 -0.400 2.040 0.895 ;
        RECT  0.000 -0.400 1.700 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 4.640 7.260 5.440 ;
        RECT  4.955 4.025 5.185 5.440 ;
        RECT  2.760 4.640 4.955 5.440 ;
        RECT  2.420 4.465 2.760 5.440 ;
        RECT  0.520 4.640 2.420 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.185 1.925 5.415 2.645 ;
        RECT  3.700 2.415 5.185 2.645 ;
        RECT  3.470 1.360 3.700 2.645 ;
        RECT  1.675 1.360 3.470 1.590 ;
        RECT  1.445 1.360 1.675 3.195 ;
        RECT  0.975 1.360 1.445 1.590 ;
        RECT  1.300 2.965 1.445 3.195 ;
    END
END AOI2BB1X4

MACRO AOI2BB1X2
    CLASS CORE ;
    FOREIGN AOI2BB1X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB1XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 1.355 4.305 3.215 ;
        RECT  2.855 1.355 4.075 1.585 ;
        RECT  3.085 2.985 4.075 3.215 ;
        RECT  2.960 2.985 3.085 3.755 ;
        RECT  2.620 2.985 2.960 3.795 ;
        RECT  2.625 1.260 2.855 1.585 ;
        RECT  2.395 0.680 2.625 1.585 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.585 1.845 3.815 2.680 ;
        RECT  2.385 1.845 3.585 2.075 ;
        RECT  2.155 1.845 2.385 2.260 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.690 2.330 1.375 2.740 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.260 0.530 1.800 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 -0.400 4.620 0.400 ;
        RECT  3.100 -0.400 3.440 0.575 ;
        RECT  1.960 -0.400 3.100 0.400 ;
        RECT  1.620 -0.400 1.960 0.895 ;
        RECT  0.520 -0.400 1.620 0.400 ;
        RECT  0.180 -0.400 0.520 0.895 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.240 4.640 4.620 5.440 ;
        RECT  3.900 3.550 4.240 5.440 ;
        RECT  1.640 4.640 3.900 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.000 4.640 1.300 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.840 2.505 3.200 2.735 ;
        RECT  1.610 1.795 1.840 3.200 ;
        RECT  1.185 1.795 1.610 2.025 ;
        RECT  0.520 2.970 1.610 3.200 ;
        RECT  0.955 0.770 1.185 2.025 ;
        RECT  0.180 2.970 0.520 3.780 ;
    END
END AOI2BB1X2

MACRO AOI2BB1X1
    CLASS CORE ;
    FOREIGN AOI2BB1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB1XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.225 3.085 3.195 ;
        RECT  2.855 1.225 2.910 4.140 ;
        RECT  2.090 1.225 2.855 1.455 ;
        RECT  2.680 2.965 2.855 4.140 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 2.795 1.965 3.195 ;
        RECT  1.315 2.795 1.960 3.220 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 1.780 1.180 2.120 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.380 0.800 2.850 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 -0.400 3.300 0.400 ;
        RECT  0.930 -0.400 1.270 0.575 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 4.640 3.300 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.000 4.640 1.300 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.430 2.105 2.620 2.465 ;
        RECT  2.200 1.875 2.430 3.755 ;
        RECT  1.695 1.875 2.200 2.105 ;
        RECT  0.180 3.525 2.200 3.755 ;
        RECT  1.465 1.305 1.695 2.105 ;
        RECT  0.450 1.305 1.465 1.535 ;
    END
END AOI2BB1X1

MACRO AOI22XL
    CLASS CORE ;
    FOREIGN AOI22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.185 3.160 3.425 ;
        RECT  2.855 1.185 2.930 1.515 ;
        RECT  2.440 3.195 2.930 3.425 ;
        RECT  1.840 1.185 2.855 1.415 ;
        RECT  2.100 3.140 2.440 3.480 ;
        RECT  1.500 1.130 1.840 1.470 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.665 0.620 2.145 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 2.350 1.530 2.725 ;
        RECT  0.800 2.380 1.190 2.725 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.625 2.400 2.680 2.740 ;
        RECT  2.080 2.360 2.625 2.740 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 1.785 2.210 2.100 ;
        RECT  1.765 1.730 2.205 2.100 ;
        RECT  1.530 1.785 1.765 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 -0.400 3.300 0.400 ;
        RECT  2.740 -0.400 3.080 0.575 ;
        RECT  0.520 -0.400 2.740 0.400 ;
        RECT  0.180 -0.400 0.520 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 4.640 3.300 5.440 ;
        RECT  0.230 4.465 0.645 5.440 ;
        RECT  0.000 4.640 0.230 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.660 4.175 3.010 4.405 ;
        RECT  1.430 3.200 1.660 4.405 ;
        RECT  0.520 3.200 1.430 3.430 ;
        RECT  0.180 3.145 0.520 3.485 ;
    END
END AOI22XL

MACRO AOI22X4
    CLASS CORE ;
    FOREIGN AOI22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI22XL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.440 1.845 8.670 4.135 ;
        RECT  8.365 1.260 8.440 2.660 ;
        RECT  7.480 3.905 8.440 4.135 ;
        RECT  8.060 1.205 8.365 2.660 ;
        RECT  0.180 1.205 8.060 1.435 ;
        RECT  7.165 3.905 7.480 4.340 ;
        RECT  7.040 4.060 7.165 4.340 ;
        RECT  4.660 4.110 7.040 4.340 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.940 1.840 3.995 2.070 ;
        RECT  3.710 1.840 3.940 2.075 ;
        RECT  0.875 1.845 3.710 2.075 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.465 2.845 2.695 ;
        RECT  2.195 2.405 2.425 2.695 ;
        RECT  0.420 2.465 2.195 2.695 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.760 1.845 6.920 2.075 ;
        RECT  4.610 1.845 4.760 2.100 ;
        RECT  4.380 1.845 4.610 2.745 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.550 2.115 7.780 2.635 ;
        RECT  5.065 2.405 7.550 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.920 -0.400 9.240 0.400 ;
        RECT  6.580 -0.400 6.920 0.915 ;
        RECT  4.360 -0.400 6.580 0.400 ;
        RECT  4.020 -0.400 4.360 0.915 ;
        RECT  1.800 -0.400 4.020 0.400 ;
        RECT  1.460 -0.400 1.800 0.915 ;
        RECT  0.000 -0.400 1.460 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 4.640 9.240 5.440 ;
        RECT  3.380 4.055 3.720 5.440 ;
        RECT  2.440 4.640 3.380 5.440 ;
        RECT  2.100 4.055 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 4.055 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.180 3.095 8.200 3.325 ;
    END
END AOI22X4

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI22XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.350 5.725 3.195 ;
        RECT  1.460 1.350 5.495 1.580 ;
        RECT  5.080 2.965 5.495 3.195 ;
        RECT  4.835 2.965 5.080 3.315 ;
        RECT  3.460 3.085 4.835 3.315 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.915 2.655 2.415 ;
        RECT  1.105 1.915 2.425 2.145 ;
        RECT  0.915 1.845 1.105 2.145 ;
        RECT  0.685 1.845 0.915 2.360 ;
        RECT  0.420 2.070 0.685 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 2.405 1.765 2.785 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.035 1.840 5.265 2.315 ;
        RECT  3.745 1.840 5.035 2.070 ;
        RECT  3.505 1.840 3.745 2.075 ;
        RECT  3.275 1.840 3.505 2.790 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.940 2.380 4.480 2.775 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.360 -0.400 5.940 0.400 ;
        RECT  5.020 -0.400 5.360 0.575 ;
        RECT  2.920 -0.400 5.020 0.400 ;
        RECT  2.580 -0.400 2.920 0.575 ;
        RECT  0.520 -0.400 2.580 0.400 ;
        RECT  0.180 -0.400 0.520 1.345 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 4.640 5.940 5.440 ;
        RECT  2.100 3.665 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 3.665 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.025 3.720 5.720 3.950 ;
        RECT  3.025 3.075 3.080 3.305 ;
        RECT  2.795 3.075 3.025 3.950 ;
        RECT  0.180 3.075 2.795 3.305 ;
    END
END AOI22X2

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI22XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.115 3.160 3.165 ;
        RECT  2.855 1.115 2.930 1.515 ;
        RECT  2.480 2.935 2.930 3.165 ;
        RECT  1.800 1.115 2.855 1.345 ;
        RECT  2.140 2.935 2.480 3.275 ;
        RECT  1.460 1.060 1.800 1.400 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.190 1.770 0.530 2.475 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.380 1.520 2.785 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 2.260 2.680 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.830 1.655 2.170 1.995 ;
        RECT  1.765 1.710 1.830 1.995 ;
        RECT  1.535 1.710 1.765 2.075 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 -0.400 3.300 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  0.520 -0.400 2.780 0.400 ;
        RECT  0.180 -0.400 0.520 1.450 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 3.300 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.780 3.585 3.120 3.925 ;
        RECT  1.840 3.695 2.780 3.925 ;
        RECT  1.500 3.635 1.840 3.975 ;
        RECT  0.520 3.690 1.500 3.920 ;
        RECT  0.180 3.050 0.520 3.920 ;
    END
END AOI22X1

MACRO AOI222XL
    CLASS CORE ;
    FOREIGN AOI222XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.135 5.065 3.095 ;
        RECT  0.180 1.135 4.835 1.365 ;
        RECT  4.760 2.635 4.835 3.095 ;
        RECT  3.965 2.865 4.760 3.095 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.385 1.270 2.885 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.520 2.370 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.525 1.725 2.075 2.100 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.595 1.820 3.145 2.200 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.170 1.845 4.520 2.540 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 1.645 3.855 2.195 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 -0.400 5.280 0.400 ;
        RECT  4.510 -0.400 4.850 0.575 ;
        RECT  1.885 -0.400 4.510 0.400 ;
        RECT  1.545 -0.400 1.885 0.905 ;
        RECT  0.000 -0.400 1.545 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 4.640 5.280 5.440 ;
        RECT  0.820 4.410 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.080 4.145 4.865 4.375 ;
        RECT  0.740 3.365 2.980 3.595 ;
    END
END AOI222XL

MACRO AOI222X4
    CLASS CORE ;
    FOREIGN AOI222X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI222XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.070 2.380 7.120 3.780 ;
        RECT  6.840 1.410 7.070 3.780 ;
        RECT  6.740 1.410 6.840 1.850 ;
        RECT  6.740 2.380 6.840 3.780 ;
        RECT  6.500 1.410 6.740 1.640 ;
        RECT  6.500 2.775 6.740 3.115 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.520 2.620 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 1.605 1.560 2.075 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 2.405 2.420 2.635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.120 3.160 2.845 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.125 2.200 4.480 2.880 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 1.670 3.820 2.335 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.480 -0.400 7.920 0.400 ;
        RECT  7.140 -0.400 7.480 0.955 ;
        RECT  6.160 -0.400 7.140 0.400 ;
        RECT  5.820 -0.400 6.160 0.955 ;
        RECT  4.740 -0.400 5.820 0.400 ;
        RECT  4.400 -0.400 4.740 0.575 ;
        RECT  2.500 -0.400 4.400 0.400 ;
        RECT  2.160 -0.400 2.500 0.575 ;
        RECT  0.680 -0.400 2.160 0.400 ;
        RECT  0.520 -0.400 0.680 0.410 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.480 4.640 7.920 5.440 ;
        RECT  7.140 4.060 7.480 5.440 ;
        RECT  6.200 4.640 7.140 5.440 ;
        RECT  5.860 3.750 6.200 5.440 ;
        RECT  1.640 4.640 5.860 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.520 4.640 1.300 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.015 2.225 6.505 2.455 ;
        RECT  5.785 1.205 6.015 2.960 ;
        RECT  5.100 1.205 5.785 1.435 ;
        RECT  5.425 2.730 5.785 2.960 ;
        RECT  4.940 2.185 5.470 2.415 ;
        RECT  5.195 2.730 5.425 3.110 ;
        RECT  4.710 1.695 4.940 3.500 ;
        RECT  2.000 4.180 4.780 4.410 ;
        RECT  4.295 1.695 4.710 1.925 ;
        RECT  3.880 3.270 4.710 3.500 ;
        RECT  4.065 1.115 4.295 1.925 ;
        RECT  3.630 1.115 4.065 1.345 ;
        RECT  3.280 0.990 3.630 1.345 ;
        RECT  1.460 0.990 3.280 1.220 ;
        RECT  0.740 3.410 2.900 3.640 ;
    END
END AOI222X4

MACRO AOI222X2
    CLASS CORE ;
    FOREIGN AOI222X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI222XL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.635 1.125 8.865 3.120 ;
        RECT  8.365 1.125 8.635 1.540 ;
        RECT  8.365 2.890 8.635 3.120 ;
        RECT  7.480 1.125 8.365 1.355 ;
        RECT  8.135 2.890 8.365 3.195 ;
        RECT  6.640 2.890 8.135 3.120 ;
        RECT  7.040 1.045 7.480 1.355 ;
        RECT  4.870 1.125 7.040 1.355 ;
        RECT  4.400 1.045 4.870 1.355 ;
        RECT  1.460 1.125 4.400 1.355 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 2.335 2.680 2.605 ;
        RECT  1.105 2.375 2.320 2.605 ;
        RECT  0.575 2.375 1.105 2.635 ;
        RECT  0.345 2.190 0.575 2.635 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.670 1.910 2.130 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 1.845 5.760 2.075 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 2.345 4.920 2.635 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.170 1.845 8.400 2.290 ;
        RECT  6.155 1.845 8.170 2.075 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.705 2.335 7.450 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.695 -0.400 9.240 0.400 ;
        RECT  8.355 -0.400 8.695 0.895 ;
        RECT  6.130 -0.400 8.355 0.400 ;
        RECT  5.790 -0.400 6.130 0.895 ;
        RECT  3.230 -0.400 5.790 0.400 ;
        RECT  2.890 -0.400 3.230 0.895 ;
        RECT  0.520 -0.400 2.890 0.400 ;
        RECT  0.180 -0.400 0.520 1.220 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 4.640 9.240 5.440 ;
        RECT  2.740 3.765 3.080 5.440 ;
        RECT  1.800 4.640 2.740 5.440 ;
        RECT  1.460 3.765 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.765 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.440 3.820 8.900 4.050 ;
        RECT  0.820 2.890 5.700 3.120 ;
    END
END AOI222X2

MACRO AOI222X1
    CLASS CORE ;
    FOREIGN AOI222X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI222XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 1.180 5.065 3.120 ;
        RECT  0.180 1.180 4.835 1.410 ;
        RECT  4.085 2.890 4.835 3.120 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.700 1.435 2.130 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.845 0.460 2.660 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 2.125 2.210 2.635 ;
        RECT  1.535 2.405 1.840 2.635 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.645 1.820 3.160 2.245 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.820 4.480 2.465 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 1.865 3.820 2.635 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.785 -0.400 5.280 0.400 ;
        RECT  4.445 -0.400 4.785 0.575 ;
        RECT  1.915 -0.400 4.445 0.400 ;
        RECT  1.575 -0.400 1.915 0.575 ;
        RECT  0.000 -0.400 1.575 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 4.640 5.280 5.440 ;
        RECT  1.460 3.790 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.890 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.165 3.820 5.065 4.050 ;
        RECT  2.665 2.875 3.145 3.105 ;
        RECT  2.435 2.875 2.665 3.430 ;
        RECT  0.820 3.200 2.435 3.430 ;
    END
END AOI222X1

MACRO AOI221XL
    CLASS CORE ;
    FOREIGN AOI221XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 0.990 4.405 3.120 ;
        RECT  4.100 0.990 4.175 1.285 ;
        RECT  3.880 2.890 4.175 3.120 ;
        RECT  2.175 0.990 4.100 1.220 ;
        RECT  1.945 0.675 2.175 1.220 ;
        RECT  1.765 0.675 1.945 0.980 ;
        RECT  1.460 0.675 1.765 0.905 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 2.405 3.745 2.635 ;
        RECT  3.390 1.820 3.620 2.635 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.315 0.520 2.100 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.360 1.340 2.820 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.565 1.570 3.085 2.075 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 1.845 1.965 2.575 ;
        RECT  1.535 1.845 1.735 2.075 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 -0.400 4.620 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  0.520 -0.400 2.780 0.400 ;
        RECT  0.180 -0.400 0.520 0.895 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 4.640 4.620 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.520 4.640 1.300 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.000 4.180 3.460 4.410 ;
        RECT  2.560 2.820 2.900 3.640 ;
        RECT  1.080 3.410 2.560 3.640 ;
        RECT  0.740 3.110 1.080 3.930 ;
    END
END AOI221XL

MACRO AOI221X4
    CLASS CORE ;
    FOREIGN AOI221X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI221XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 1.260 6.460 2.660 ;
        RECT  6.080 1.260 6.310 4.050 ;
        RECT  5.900 1.260 6.080 1.490 ;
        RECT  5.960 2.770 6.080 4.050 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 1.565 3.745 2.075 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.940 0.520 2.655 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.510 1.220 3.195 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.655 2.380 3.085 2.635 ;
        RECT  2.425 2.110 2.655 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 1.820 1.940 2.455 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.920 -0.400 7.260 0.400 ;
        RECT  6.690 -0.400 6.920 1.580 ;
        RECT  5.520 -0.400 6.690 0.400 ;
        RECT  5.180 -0.400 5.520 0.895 ;
        RECT  3.120 -0.400 5.180 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  0.520 -0.400 2.780 0.400 ;
        RECT  0.180 -0.400 0.520 1.285 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.020 4.640 7.260 5.440 ;
        RECT  6.680 3.150 7.020 5.440 ;
        RECT  5.580 4.640 6.680 5.440 ;
        RECT  5.240 3.150 5.580 5.440 ;
        RECT  1.640 4.640 5.240 5.440 ;
        RECT  1.300 4.465 1.640 5.440 ;
        RECT  0.520 4.640 1.300 5.440 ;
        RECT  0.180 4.465 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.070 2.135 5.710 2.365 ;
        RECT  4.860 1.450 5.070 2.705 ;
        RECT  4.840 1.450 4.860 4.100 ;
        RECT  4.740 1.450 4.840 1.680 ;
        RECT  4.630 2.475 4.840 4.100 ;
        RECT  4.510 1.150 4.740 1.680 ;
        RECT  4.520 3.760 4.630 4.100 ;
        RECT  4.280 1.965 4.610 2.195 ;
        RECT  4.050 0.990 4.280 3.400 ;
        RECT  2.415 0.990 4.050 1.220 ;
        RECT  3.935 3.035 4.050 3.400 ;
        RECT  0.740 3.495 2.900 3.725 ;
        RECT  2.185 0.990 2.415 1.285 ;
        RECT  1.460 1.055 2.185 1.285 ;
    END
END AOI221X4

MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI221XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.310 7.045 3.510 ;
        RECT  5.495 1.310 6.815 1.540 ;
        RECT  6.640 3.170 6.815 3.510 ;
        RECT  5.245 1.260 5.495 1.540 ;
        RECT  5.015 0.945 5.245 1.540 ;
        RECT  1.460 0.945 5.015 1.175 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.330 1.845 6.560 2.280 ;
        RECT  5.495 1.845 6.330 2.075 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 2.070 2.680 2.345 ;
        RECT  2.120 1.820 2.500 2.345 ;
        RECT  0.290 2.115 2.120 2.345 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.575 1.560 1.805 ;
        RECT  0.800 1.285 1.180 1.805 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 2.500 5.930 2.730 ;
        RECT  3.515 2.405 3.745 2.730 ;
        RECT  3.460 2.500 3.515 2.730 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.665 4.650 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.170 -0.400 7.920 0.400 ;
        RECT  5.830 -0.400 6.170 0.895 ;
        RECT  3.280 -0.400 5.830 0.400 ;
        RECT  2.940 -0.400 3.280 0.575 ;
        RECT  0.520 -0.400 2.940 0.400 ;
        RECT  0.180 -0.400 0.520 0.895 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 4.640 7.920 5.440 ;
        RECT  2.740 3.730 3.080 5.440 ;
        RECT  1.800 4.640 2.740 5.440 ;
        RECT  1.460 3.730 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.730 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.440 4.040 7.620 4.270 ;
        RECT  3.560 3.225 5.700 3.455 ;
        RECT  3.330 2.970 3.560 3.455 ;
        RECT  0.820 2.970 3.330 3.200 ;
    END
END AOI221X2

MACRO AOI221X1
    CLASS CORE ;
    FOREIGN AOI221X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI221XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 1.080 4.405 3.195 ;
        RECT  2.500 1.080 4.175 1.310 ;
        RECT  4.140 2.635 4.175 3.165 ;
        RECT  2.475 0.955 2.500 1.310 ;
        RECT  2.245 0.795 2.475 1.310 ;
        RECT  1.460 0.795 2.245 1.025 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.710 2.405 3.745 2.635 ;
        RECT  3.480 1.650 3.710 2.635 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.175 1.285 0.520 1.935 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.185 1.350 2.660 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.590 3.085 2.075 ;
        RECT  2.370 1.590 2.855 1.820 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.535 1.285 1.990 1.810 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 -0.400 4.620 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  0.520 -0.400 2.780 0.400 ;
        RECT  0.180 -0.400 0.520 1.025 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 4.640 4.620 5.440 ;
        RECT  1.460 3.785 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 3.785 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.165 3.620 3.785 3.850 ;
        RECT  0.820 2.895 3.145 3.125 ;
    END
END AOI221X1

MACRO AOI21XL
    CLASS CORE ;
    FOREIGN AOI21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.390 1.240 2.425 2.635 ;
        RECT  2.195 1.240 2.390 3.485 ;
        RECT  1.460 1.240 2.195 1.470 ;
        RECT  2.160 2.405 2.195 3.485 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.365 1.725 1.935 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.170 1.750 0.520 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.380 1.430 2.780 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 -0.400 2.640 0.400 ;
        RECT  2.020 -0.400 2.360 0.575 ;
        RECT  0.520 -0.400 2.020 0.400 ;
        RECT  0.180 -0.400 0.520 1.455 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 4.640 2.640 5.440 ;
        RECT  0.840 4.465 1.180 5.440 ;
        RECT  0.000 4.640 0.840 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.640 4.180 1.880 4.410 ;
        RECT  1.410 4.000 1.640 4.410 ;
        RECT  0.465 4.000 1.410 4.230 ;
        RECT  0.235 3.145 0.465 4.230 ;
    END
END AOI21XL

MACRO AOI21X4
    CLASS CORE ;
    FOREIGN AOI21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI21XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.115 3.765 6.280 4.105 ;
        RECT  5.940 2.430 6.115 4.105 ;
        RECT  5.885 2.430 5.940 4.050 ;
        RECT  5.800 2.430 5.885 2.660 ;
        RECT  5.000 3.820 5.885 4.050 ;
        RECT  5.420 1.260 5.800 2.660 ;
        RECT  4.835 1.415 5.420 1.645 ;
        RECT  4.660 3.765 5.000 4.105 ;
        RECT  4.430 1.150 4.835 1.645 ;
        RECT  0.180 1.150 4.430 1.380 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 2.085 5.140 2.665 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.915 1.900 4.025 2.240 ;
        RECT  3.685 1.645 3.915 2.240 ;
        RECT  2.425 1.645 3.685 1.875 ;
        RECT  1.805 1.645 2.425 2.075 ;
        RECT  1.520 1.645 1.805 2.130 ;
        RECT  1.465 1.790 1.520 2.130 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 2.405 3.085 2.635 ;
        RECT  2.730 2.225 2.960 2.635 ;
        RECT  0.800 2.395 2.730 2.625 ;
        RECT  0.760 2.380 0.800 2.625 ;
        RECT  0.530 1.970 0.760 2.625 ;
        RECT  0.420 1.970 0.530 2.410 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.685 -0.400 6.600 0.400 ;
        RECT  5.345 -0.400 5.685 0.575 ;
        RECT  4.365 -0.400 5.345 0.400 ;
        RECT  4.025 -0.400 4.365 0.895 ;
        RECT  1.805 -0.400 4.025 0.400 ;
        RECT  1.465 -0.400 1.805 0.895 ;
        RECT  0.000 -0.400 1.465 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 4.640 6.600 5.440 ;
        RECT  3.380 3.890 3.720 5.440 ;
        RECT  2.440 4.640 3.380 5.440 ;
        RECT  2.100 3.890 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 3.890 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.180 2.930 5.640 3.160 ;
    END
END AOI21X4

MACRO AOI21X2
    CLASS CORE ;
    FOREIGN AOI21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI21XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.660 1.450 3.890 3.315 ;
        RECT  3.080 1.450 3.660 1.680 ;
        RECT  3.515 2.965 3.660 3.315 ;
        RECT  3.460 3.085 3.515 3.315 ;
        RECT  2.740 1.125 3.080 1.680 ;
        RECT  1.065 1.450 2.740 1.680 ;
        RECT  0.835 1.235 1.065 1.680 ;
        RECT  0.520 1.235 0.835 1.465 ;
        RECT  0.180 1.125 0.520 1.465 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 2.035 3.325 2.635 ;
        RECT  2.855 2.405 2.950 2.635 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.500 1.840 2.810 ;
        RECT  0.875 2.405 1.105 2.810 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 1.920 2.710 2.150 ;
        RECT  0.140 1.820 0.520 2.225 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.845 -0.400 4.620 0.400 ;
        RECT  3.505 -0.400 3.845 0.575 ;
        RECT  1.800 -0.400 3.505 0.400 ;
        RECT  1.460 -0.400 1.800 1.220 ;
        RECT  0.000 -0.400 1.460 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 4.640 4.620 5.440 ;
        RECT  2.100 3.665 2.440 5.440 ;
        RECT  1.160 4.640 2.100 5.440 ;
        RECT  0.820 3.665 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.100 3.665 4.440 4.005 ;
        RECT  3.095 3.665 4.100 3.895 ;
        RECT  2.865 3.075 3.095 3.895 ;
        RECT  0.180 3.075 2.865 3.305 ;
    END
END AOI21X2

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI21XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.275 1.350 2.505 3.950 ;
        RECT  1.800 1.350 2.275 1.580 ;
        RECT  2.195 2.965 2.275 3.950 ;
        RECT  2.100 3.610 2.195 3.950 ;
        RECT  1.460 1.240 1.800 1.580 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 1.845 2.045 2.635 ;
        RECT  1.535 1.845 1.800 2.075 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.065 0.530 2.585 ;
        RECT  0.190 1.820 0.520 2.585 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.385 1.430 2.615 ;
        RECT  0.875 1.285 1.105 2.615 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 -0.400 2.640 0.400 ;
        RECT  2.020 -0.400 2.360 0.575 ;
        RECT  0.520 -0.400 2.020 0.400 ;
        RECT  0.180 -0.400 0.520 1.465 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 4.640 2.640 5.440 ;
        RECT  0.820 3.515 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.180 2.925 1.800 3.155 ;
    END
END AOI21X1

MACRO AOI211XL
    CLASS CORE ;
    FOREIGN AOI211XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.150 3.160 3.195 ;
        RECT  1.460 1.150 2.930 1.380 ;
        RECT  2.780 2.965 2.930 3.195 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.510 2.330 2.125 2.710 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.470 1.820 2.700 2.485 ;
        RECT  2.115 1.820 2.470 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.955 0.520 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.650 1.375 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 -0.400 3.300 0.400 ;
        RECT  2.120 -0.400 2.460 0.575 ;
        RECT  0.520 -0.400 2.120 0.400 ;
        RECT  0.180 -0.400 0.520 1.240 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 4.640 3.300 5.440 ;
        RECT  0.740 4.465 1.080 5.440 ;
        RECT  0.000 4.640 0.740 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.180 2.955 1.840 3.185 ;
    END
END AOI211XL

MACRO AOI211X4
    CLASS CORE ;
    FOREIGN AOI211X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI211XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.140 0.760 5.325 1.585 ;
        RECT  5.140 2.740 5.195 3.080 ;
        RECT  5.095 0.760 5.140 3.080 ;
        RECT  4.855 1.260 5.095 3.080 ;
        RECT  4.760 1.260 4.855 2.660 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 2.380 2.070 2.710 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.415 3.160 3.220 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.215 1.285 0.495 2.100 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.775 1.440 2.100 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.100 -0.400 6.600 0.400 ;
        RECT  5.760 -0.400 6.100 1.420 ;
        RECT  4.660 -0.400 5.760 0.400 ;
        RECT  4.320 -0.400 4.660 0.895 ;
        RECT  2.340 -0.400 4.320 0.400 ;
        RECT  2.000 -0.400 2.340 0.575 ;
        RECT  0.520 -0.400 2.000 0.400 ;
        RECT  0.180 -0.400 0.520 0.895 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 4.640 6.600 5.440 ;
        RECT  5.495 4.010 5.835 5.440 ;
        RECT  4.555 4.640 5.495 5.440 ;
        RECT  4.215 3.815 4.555 5.440 ;
        RECT  1.085 4.640 4.215 5.440 ;
        RECT  0.745 4.465 1.085 5.440 ;
        RECT  0.000 4.640 0.745 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.600 2.180 5.830 3.580 ;
        RECT  4.315 3.350 5.600 3.580 ;
        RECT  4.085 1.135 4.315 3.580 ;
        RECT  3.885 1.135 4.085 1.365 ;
        RECT  3.835 3.055 4.085 3.580 ;
        RECT  3.655 0.880 3.885 1.365 ;
        RECT  3.295 1.735 3.850 1.965 ;
        RECT  3.495 3.055 3.835 3.875 ;
        RECT  3.065 1.130 3.295 1.965 ;
        RECT  2.530 3.465 3.130 3.695 ;
        RECT  1.500 1.130 3.065 1.360 ;
        RECT  2.530 1.735 3.065 1.965 ;
        RECT  2.300 1.735 2.530 3.695 ;
        RECT  0.180 3.235 1.850 3.465 ;
    END
END AOI211X4

MACRO AOI211X2
    CLASS CORE ;
    FOREIGN AOI211X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI211XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 1.045 5.690 3.195 ;
        RECT  5.250 1.045 5.460 1.275 ;
        RECT  4.370 2.965 5.460 3.195 ;
        RECT  4.910 0.935 5.250 1.275 ;
        RECT  3.640 0.990 4.910 1.220 ;
        RECT  4.085 2.965 4.370 3.390 ;
        RECT  4.030 3.050 4.085 3.390 ;
        RECT  2.830 0.935 3.640 1.275 ;
        RECT  2.780 0.935 2.830 1.220 ;
        RECT  0.530 0.990 2.780 1.220 ;
        RECT  0.190 0.935 0.530 1.275 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.995 1.535 5.225 2.265 ;
        RECT  4.760 1.535 4.995 1.845 ;
        RECT  3.360 1.535 4.760 1.765 ;
        RECT  3.130 1.535 3.360 2.635 ;
        RECT  2.855 2.310 3.130 2.635 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 2.310 4.480 2.710 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 2.265 1.480 2.635 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 2.075 2.285 2.610 ;
        RECT  2.000 1.675 2.230 2.610 ;
        RECT  0.770 1.675 2.000 1.905 ;
        RECT  1.945 2.270 2.000 2.610 ;
        RECT  0.445 1.620 0.770 1.960 ;
        RECT  0.430 1.620 0.445 2.075 ;
        RECT  0.215 1.675 0.430 2.075 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.485 -0.400 5.940 0.400 ;
        RECT  4.145 -0.400 4.485 0.575 ;
        RECT  1.850 -0.400 4.145 0.400 ;
        RECT  1.510 -0.400 1.850 0.575 ;
        RECT  0.000 -0.400 1.510 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.445 4.640 5.940 5.440 ;
        RECT  2.105 3.820 2.445 5.440 ;
        RECT  1.165 4.640 2.105 5.440 ;
        RECT  0.825 3.820 1.165 5.440 ;
        RECT  0.000 4.640 0.825 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.310 3.700 5.650 4.040 ;
        RECT  3.480 3.755 5.310 3.985 ;
        RECT  3.250 2.890 3.480 3.985 ;
        RECT  0.185 2.890 3.250 3.120 ;
    END
END AOI211X2

MACRO AOI211X1
    CLASS CORE ;
    FOREIGN AOI211X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI211XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 1.095 3.180 3.195 ;
        RECT  3.010 1.095 3.080 4.095 ;
        RECT  2.950 0.805 3.010 4.095 ;
        RECT  2.780 0.805 2.950 1.435 ;
        RECT  2.740 2.775 2.950 4.095 ;
        RECT  1.835 0.805 2.780 1.035 ;
        RECT  1.605 0.805 1.835 1.380 ;
        RECT  1.460 1.150 1.605 1.380 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.165 2.045 2.660 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 1.830 2.720 2.250 ;
        RECT  2.490 1.830 2.510 3.195 ;
        RECT  2.280 2.020 2.490 3.195 ;
        RECT  2.195 2.965 2.280 3.195 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.200 0.645 2.710 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.680 1.430 1.910 ;
        RECT  0.875 1.285 1.180 1.910 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.345 -0.400 3.300 0.400 ;
        RECT  2.005 -0.400 2.345 0.575 ;
        RECT  0.520 -0.400 2.005 0.400 ;
        RECT  0.180 -0.400 0.520 1.155 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 4.640 3.300 5.440 ;
        RECT  0.820 3.755 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.180 3.115 1.800 3.345 ;
    END
END AOI211X1

MACRO AND4XL
    CLASS CORE ;
    FOREIGN AND4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.705 3.190 3.820 3.780 ;
        RECT  3.475 1.015 3.705 3.780 ;
        RECT  3.420 3.190 3.475 3.780 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.540 2.405 3.105 2.890 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.135 1.840 2.890 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.135 1.180 2.890 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.545 0.520 3.220 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.000 -0.400 3.960 0.400 ;
        RECT  2.660 -0.400 3.000 0.575 ;
        RECT  0.000 -0.400 2.660 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.100 4.640 3.960 5.440 ;
        RECT  0.930 4.465 3.100 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.300 1.540 3.225 1.910 ;
        RECT  2.260 0.975 2.300 3.460 ;
        RECT  2.070 0.975 2.260 3.725 ;
        RECT  0.520 0.975 2.070 1.205 ;
        RECT  1.920 3.155 2.070 3.725 ;
        RECT  0.520 3.495 1.920 3.725 ;
        RECT  0.180 0.975 0.520 1.315 ;
    END
END AND4XL

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND4XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.385 2.380 6.460 3.780 ;
        RECT  6.155 1.495 6.385 3.780 ;
        RECT  6.085 1.390 6.155 3.780 ;
        RECT  6.080 1.390 6.085 1.845 ;
        RECT  6.080 2.380 6.085 3.780 ;
        RECT  5.700 1.390 6.080 1.730 ;
        RECT  5.560 3.425 6.080 3.780 ;
        RECT  5.220 3.425 5.560 4.365 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.845 4.950 2.075 ;
        RECT  4.590 1.845 4.820 2.730 ;
        RECT  4.405 2.380 4.590 2.730 ;
        RECT  4.275 2.500 4.405 2.730 ;
        RECT  4.045 2.500 4.275 3.730 ;
        RECT  0.525 3.500 4.045 3.730 ;
        RECT  0.525 2.690 0.530 3.220 ;
        RECT  0.295 2.690 0.525 3.730 ;
        RECT  0.140 2.690 0.295 3.220 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.585 1.590 3.815 3.030 ;
        RECT  3.440 1.590 3.585 1.845 ;
        RECT  1.250 1.590 3.440 1.820 ;
        RECT  1.250 2.265 1.320 2.670 ;
        RECT  1.020 1.590 1.250 2.670 ;
        RECT  0.800 2.070 1.020 2.670 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 2.055 3.160 2.640 ;
        RECT  1.670 2.055 2.780 2.285 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.625 2.500 3.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.760 -0.400 7.260 0.400 ;
        RECT  6.420 -0.400 6.760 0.950 ;
        RECT  5.320 -0.400 6.420 0.400 ;
        RECT  4.980 -0.400 5.320 1.115 ;
        RECT  0.520 -0.400 4.980 0.400 ;
        RECT  0.180 -0.400 0.520 1.465 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.355 4.640 7.260 5.440 ;
        RECT  5.965 4.465 6.355 5.440 ;
        RECT  4.445 4.640 5.965 5.440 ;
        RECT  4.105 4.465 4.445 5.440 ;
        RECT  2.840 4.640 4.105 5.440 ;
        RECT  2.500 4.465 2.840 5.440 ;
        RECT  1.300 4.640 2.500 5.440 ;
        RECT  0.910 4.465 1.300 5.440 ;
        RECT  0.000 4.640 0.910 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.470 2.130 5.715 2.470 ;
        RECT  5.240 1.380 5.470 3.195 ;
        RECT  4.455 1.380 5.240 1.610 ;
        RECT  4.740 2.965 5.240 3.195 ;
        RECT  4.510 2.965 4.740 4.195 ;
        RECT  3.625 3.965 4.510 4.195 ;
        RECT  4.225 1.065 4.455 1.610 ;
        RECT  2.920 1.065 4.225 1.295 ;
        RECT  3.285 3.965 3.625 4.365 ;
        RECT  2.080 3.965 3.285 4.195 ;
        RECT  2.580 1.010 2.920 1.350 ;
        RECT  1.740 3.965 2.080 4.365 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.775 2.940 3.820 3.220 ;
        RECT  3.710 1.505 3.775 3.220 ;
        RECT  3.545 0.835 3.710 4.050 ;
        RECT  3.480 0.835 3.545 1.735 ;
        RECT  3.480 2.720 3.545 4.050 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.500 2.200 2.640 2.545 ;
        RECT  2.195 1.845 2.500 2.545 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.720 2.440 1.950 3.195 ;
        RECT  1.535 2.965 1.720 3.195 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 2.255 1.290 2.715 ;
        RECT  0.800 2.255 1.005 2.710 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.670 0.565 2.335 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 -0.400 3.960 0.400 ;
        RECT  2.595 -0.400 2.935 0.575 ;
        RECT  0.000 -0.400 2.595 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.015 4.640 3.960 5.440 ;
        RECT  2.605 4.405 3.015 5.440 ;
        RECT  1.850 4.640 2.605 5.440 ;
        RECT  1.510 4.465 1.850 5.440 ;
        RECT  0.570 4.640 1.510 5.440 ;
        RECT  0.175 4.465 0.570 5.440 ;
        RECT  0.000 4.640 0.175 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.200 1.985 3.310 2.335 ;
        RECT  2.970 0.885 3.200 3.735 ;
        RECT  0.560 0.885 2.970 1.115 ;
        RECT  0.750 3.505 2.970 3.735 ;
        RECT  0.275 0.885 0.560 1.440 ;
        RECT  0.220 1.050 0.275 1.440 ;
    END
END AND4X2

MACRO AND4X1
    CLASS CORE ;
    FOREIGN AND4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 3.195 3.820 3.800 ;
        RECT  3.530 1.025 3.760 3.800 ;
        RECT  3.420 1.025 3.530 1.365 ;
        RECT  3.440 3.195 3.530 3.800 ;
        RECT  3.420 3.360 3.440 3.800 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.530 2.405 3.085 2.925 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.410 2.380 1.840 2.925 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 1.675 1.180 2.290 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.585 0.530 3.260 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.000 -0.400 3.960 0.400 ;
        RECT  2.660 -0.400 3.000 0.575 ;
        RECT  0.000 -0.400 2.660 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.100 4.640 3.960 5.440 ;
        RECT  0.930 4.465 3.100 5.440 ;
        RECT  0.000 4.640 0.930 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.160 1.685 3.270 2.025 ;
        RECT  2.930 0.935 3.160 2.025 ;
        RECT  0.520 0.935 2.930 1.165 ;
        RECT  2.300 1.740 2.930 1.970 ;
        RECT  2.260 1.740 2.300 3.460 ;
        RECT  2.070 1.740 2.260 3.725 ;
        RECT  1.920 3.155 2.070 3.725 ;
        RECT  0.520 3.495 1.920 3.725 ;
        RECT  0.180 0.935 0.520 1.275 ;
    END
END AND4X1

MACRO AND3XL
    CLASS CORE ;
    FOREIGN AND3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.150 3.495 3.160 4.240 ;
        RECT  2.920 1.150 3.150 4.240 ;
        RECT  2.780 1.150 2.920 1.490 ;
        RECT  2.740 3.495 2.920 4.240 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 1.715 1.975 2.145 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.630 2.845 1.135 3.300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.790 0.580 2.300 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 -0.400 3.300 0.400 ;
        RECT  2.000 -0.400 2.340 0.575 ;
        RECT  0.000 -0.400 2.000 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.465 4.640 3.300 5.440 ;
        RECT  2.465 2.620 2.690 3.125 ;
        RECT  2.235 2.620 2.465 5.440 ;
        RECT  1.340 4.640 2.235 5.440 ;
        RECT  1.335 4.465 1.340 5.440 ;
        RECT  1.010 4.410 1.335 5.440 ;
        RECT  1.000 4.465 1.010 5.440 ;
        RECT  0.000 4.640 1.000 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.550 1.750 2.690 2.100 ;
        RECT  2.320 1.125 2.550 2.100 ;
        RECT  1.055 1.125 2.320 1.355 ;
        RECT  1.520 2.380 1.750 4.180 ;
        RECT  1.465 2.380 1.520 3.125 ;
        RECT  0.540 3.950 1.520 4.180 ;
        RECT  1.055 2.380 1.465 2.610 ;
        RECT  0.825 1.125 1.055 2.610 ;
        RECT  0.520 1.125 0.825 1.355 ;
        RECT  0.200 3.950 0.540 4.355 ;
        RECT  0.180 1.070 0.520 1.410 ;
    END
END AND3XL

MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND3XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.820 3.820 3.220 ;
        RECT  3.440 1.690 3.745 3.220 ;
        RECT  2.985 1.690 3.440 1.920 ;
        RECT  2.850 2.800 3.440 3.155 ;
        RECT  2.755 1.375 2.985 1.920 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.835 1.820 2.065 2.420 ;
        RECT  1.460 1.820 1.835 2.100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.350 1.485 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.820 0.570 2.425 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 -0.400 3.960 0.400 ;
        RECT  3.440 -0.400 3.780 0.575 ;
        RECT  2.390 -0.400 3.440 0.400 ;
        RECT  2.050 -0.400 2.390 1.030 ;
        RECT  0.000 -0.400 2.050 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 4.640 3.960 5.440 ;
        RECT  3.440 3.855 3.780 5.440 ;
        RECT  2.460 4.640 3.440 5.440 ;
        RECT  2.120 3.750 2.460 5.440 ;
        RECT  1.160 4.640 2.120 5.440 ;
        RECT  0.820 3.750 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.525 2.295 3.065 2.525 ;
        RECT  2.295 1.330 2.525 3.370 ;
        RECT  1.605 1.330 2.295 1.560 ;
        RECT  0.180 3.140 2.295 3.370 ;
        RECT  1.375 1.135 1.605 1.560 ;
        RECT  0.535 1.135 1.375 1.365 ;
        RECT  0.195 1.080 0.535 1.420 ;
    END
END AND3X4

MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND3XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 1.330 3.100 3.195 ;
        RECT  2.870 0.790 2.960 3.195 ;
        RECT  2.620 0.790 2.870 1.610 ;
        RECT  2.815 2.740 2.870 3.195 ;
        RECT  2.760 2.740 2.815 3.080 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.870 2.520 1.980 2.895 ;
        RECT  1.640 1.820 1.870 2.895 ;
        RECT  1.460 1.820 1.640 2.100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.025 2.370 1.255 2.895 ;
        RECT  0.800 2.380 1.025 2.895 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.465 0.570 2.805 ;
        RECT  0.140 2.465 0.520 3.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 -0.400 3.300 0.400 ;
        RECT  1.860 -0.400 2.200 0.575 ;
        RECT  0.000 -0.400 1.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 4.640 3.300 5.440 ;
        RECT  2.000 4.410 2.340 5.440 ;
        RECT  0.000 4.640 2.000 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.475 2.050 2.640 2.450 ;
        RECT  2.390 2.050 2.475 3.480 ;
        RECT  2.245 1.360 2.390 3.480 ;
        RECT  2.160 1.360 2.245 2.280 ;
        RECT  1.120 3.250 2.245 3.480 ;
        RECT  0.520 1.360 2.160 1.590 ;
        RECT  0.890 3.250 1.120 4.235 ;
        RECT  0.520 4.005 0.890 4.235 ;
        RECT  0.180 1.250 0.520 1.590 ;
        RECT  0.175 4.005 0.520 4.405 ;
    END
END AND3X2

MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND3XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 1.150 3.150 4.155 ;
        RECT  2.690 1.150 2.920 1.490 ;
        RECT  2.780 3.480 2.920 4.155 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 1.715 1.975 2.145 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.675 2.845 1.180 3.300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.790 0.580 2.300 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 -0.400 3.300 0.400 ;
        RECT  2.000 -0.400 2.340 0.575 ;
        RECT  0.000 -0.400 2.000 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 4.640 3.300 5.440 ;
        RECT  2.545 2.755 2.690 3.095 ;
        RECT  2.315 2.755 2.545 5.440 ;
        RECT  1.320 4.640 2.315 5.440 ;
        RECT  1.315 4.465 1.320 5.440 ;
        RECT  0.990 4.410 1.315 5.440 ;
        RECT  0.980 4.465 0.990 5.440 ;
        RECT  0.000 4.640 0.980 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.435 1.750 2.690 2.115 ;
        RECT  2.205 1.190 2.435 2.115 ;
        RECT  1.055 1.190 2.205 1.420 ;
        RECT  1.695 2.380 1.750 3.125 ;
        RECT  1.465 2.380 1.695 4.180 ;
        RECT  1.055 2.380 1.465 2.610 ;
        RECT  0.520 3.950 1.465 4.180 ;
        RECT  0.825 1.190 1.055 2.610 ;
        RECT  0.520 1.190 0.825 1.420 ;
        RECT  0.180 1.080 0.520 1.420 ;
        RECT  0.180 3.950 0.520 4.360 ;
    END
END AND3X1

MACRO AND2XL
    CLASS CORE ;
    FOREIGN AND2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 2.380 2.500 2.660 ;
        RECT  2.125 1.445 2.355 3.550 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 2.370 1.205 2.950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 1.820 0.565 2.315 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 -0.400 2.640 0.400 ;
        RECT  1.450 -0.400 1.790 0.575 ;
        RECT  0.000 -0.400 1.450 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.400 4.640 2.640 5.440 ;
        RECT  0.460 4.465 1.400 5.440 ;
        RECT  0.000 4.640 0.460 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.660 0.820 1.890 3.475 ;
        RECT  0.520 0.820 1.660 1.050 ;
        RECT  0.800 3.245 1.660 3.475 ;
        RECT  0.460 3.190 0.800 3.530 ;
        RECT  0.180 0.765 0.520 1.105 ;
    END
END AND2XL

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 1.820 3.160 3.220 ;
        RECT  2.875 1.390 3.155 3.350 ;
        RECT  2.780 1.370 2.875 3.350 ;
        RECT  2.170 1.370 2.780 1.820 ;
        RECT  2.125 3.010 2.780 3.350 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.980 1.375 2.360 ;
        RECT  1.145 1.980 1.180 3.300 ;
        RECT  0.950 2.130 1.145 3.300 ;
        RECT  0.800 2.635 0.950 3.300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.025 0.530 2.410 ;
        RECT  0.140 2.025 0.520 2.770 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 -0.400 3.300 0.400 ;
        RECT  2.770 -0.400 3.110 1.085 ;
        RECT  1.760 -0.400 2.770 0.400 ;
        RECT  1.420 -0.400 1.760 0.575 ;
        RECT  0.000 -0.400 1.420 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.110 4.640 3.300 5.440 ;
        RECT  2.770 3.775 3.110 5.440 ;
        RECT  1.785 4.640 2.770 5.440 ;
        RECT  1.445 4.465 1.785 5.440 ;
        RECT  0.535 4.640 1.445 5.440 ;
        RECT  0.170 4.465 0.535 5.440 ;
        RECT  0.000 4.640 0.170 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.845 2.090 2.430 2.430 ;
        RECT  1.645 1.485 1.845 2.820 ;
        RECT  1.615 1.485 1.645 3.820 ;
        RECT  0.520 1.485 1.615 1.715 ;
        RECT  1.415 2.590 1.615 3.820 ;
        RECT  0.740 3.590 1.415 3.820 ;
        RECT  0.180 1.440 0.520 1.780 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND2XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.420 0.955 2.465 3.220 ;
        RECT  2.235 0.820 2.420 4.210 ;
        RECT  2.195 0.820 2.235 1.845 ;
        RECT  2.080 2.890 2.235 4.210 ;
        RECT  2.080 0.820 2.195 1.640 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 3.500 1.360 3.925 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 2.115 0.760 2.455 ;
        RECT  0.140 2.115 0.520 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.660 -0.400 2.640 0.400 ;
        RECT  1.320 -0.400 1.660 0.575 ;
        RECT  0.000 -0.400 1.320 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.570 4.640 2.640 5.440 ;
        RECT  0.180 4.465 0.570 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.225 2.150 1.965 2.495 ;
        RECT  0.995 1.460 1.225 3.095 ;
        RECT  0.520 1.460 0.995 1.690 ;
        RECT  0.815 2.745 0.995 3.095 ;
        RECT  0.180 1.350 0.520 1.690 ;
    END
END AND2X2

MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND2XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 2.380 2.500 2.660 ;
        RECT  2.355 1.345 2.410 1.845 ;
        RECT  2.355 3.075 2.410 3.895 ;
        RECT  2.125 1.345 2.355 3.895 ;
        RECT  2.120 1.345 2.125 1.845 ;
        RECT  2.070 3.075 2.125 3.895 ;
        RECT  2.070 1.345 2.120 1.685 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 2.315 1.215 2.895 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.150 1.820 0.565 2.315 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 -0.400 2.640 0.400 ;
        RECT  1.450 -0.400 1.790 0.575 ;
        RECT  0.000 -0.400 1.450 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.755 4.640 2.640 5.440 ;
        RECT  1.310 4.465 1.755 5.440 ;
        RECT  0.790 4.640 1.310 5.440 ;
        RECT  0.450 4.465 0.790 5.440 ;
        RECT  0.000 4.640 0.450 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.835 1.935 1.885 2.355 ;
        RECT  1.605 0.820 1.835 3.475 ;
        RECT  0.520 0.820 1.605 1.050 ;
        RECT  1.595 1.935 1.605 2.355 ;
        RECT  0.790 3.245 1.605 3.475 ;
        RECT  0.450 3.190 0.790 3.530 ;
        RECT  0.180 0.765 0.520 1.105 ;
    END
END AND2X1

MACRO ADDHXL
    CLASS CORE ;
    FOREIGN ADDHXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.355 2.965 4.405 3.205 ;
        RECT  4.125 1.625 4.355 3.205 ;
        RECT  3.490 1.625 4.125 1.855 ;
        RECT  3.410 2.975 4.125 3.205 ;
        RECT  3.260 1.095 3.490 1.855 ;
        RECT  3.180 2.975 3.410 3.685 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.025 1.845 7.045 2.075 ;
        RECT  6.795 0.630 7.025 3.845 ;
        RECT  6.500 3.615 6.795 3.845 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 3.930 5.745 4.160 ;
        RECT  3.605 2.135 3.835 2.740 ;
        RECT  2.950 2.510 3.605 2.740 ;
        RECT  2.720 2.510 2.950 4.160 ;
        RECT  2.120 2.865 2.720 3.220 ;
        RECT  1.775 2.865 2.120 3.095 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 2.310 5.800 2.730 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.360 -0.400 7.260 0.400 ;
        RECT  6.020 -0.400 6.360 0.970 ;
        RECT  5.065 -0.400 6.020 0.400 ;
        RECT  4.725 -0.400 5.065 0.575 ;
        RECT  1.280 -0.400 4.725 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.275 4.640 7.260 5.440 ;
        RECT  5.935 4.465 6.275 5.440 ;
        RECT  4.745 4.640 5.935 5.440 ;
        RECT  4.405 4.465 4.745 5.440 ;
        RECT  1.280 4.640 4.405 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.300 2.810 6.540 3.215 ;
        RECT  6.070 1.390 6.300 3.215 ;
        RECT  5.885 1.390 6.070 1.620 ;
        RECT  5.450 2.985 6.070 3.215 ;
        RECT  5.220 2.985 5.450 3.685 ;
        RECT  4.710 1.155 4.940 3.685 ;
        RECT  4.210 1.155 4.710 1.385 ;
        RECT  3.845 3.455 4.710 3.685 ;
        RECT  3.980 0.630 4.210 1.385 ;
        RECT  2.995 0.630 3.980 0.860 ;
        RECT  2.765 0.630 2.995 2.135 ;
        RECT  1.390 1.905 2.765 2.135 ;
        RECT  2.300 0.635 2.530 1.035 ;
        RECT  2.255 3.580 2.485 4.235 ;
        RECT  0.925 1.265 2.425 1.495 ;
        RECT  0.465 0.805 2.300 1.035 ;
        RECT  0.465 4.005 2.255 4.235 ;
        RECT  1.535 3.545 1.840 3.775 ;
        RECT  1.305 2.985 1.535 3.775 ;
        RECT  1.160 1.905 1.390 2.670 ;
        RECT  0.925 2.985 1.305 3.215 ;
        RECT  0.695 1.265 0.925 3.215 ;
        RECT  0.235 0.805 0.465 4.235 ;
    END
END ADDHXL

MACRO ADDHX4
    CLASS CORE ;
    FOREIGN ADDHX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDHXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.340 0.665 10.650 1.005 ;
        RECT  8.135 0.665 10.340 0.895 ;
        RECT  5.725 2.985 10.245 3.215 ;
        RECT  7.905 0.665 8.135 1.645 ;
        RECT  7.705 1.260 7.905 1.645 ;
        RECT  5.800 1.415 7.705 1.645 ;
        RECT  5.725 1.260 5.800 2.660 ;
        RECT  5.495 1.260 5.725 3.215 ;
        RECT  5.420 1.260 5.495 2.660 ;
        RECT  4.780 2.985 5.495 3.215 ;
        RECT  5.220 1.315 5.420 1.700 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.530 2.380 17.680 3.780 ;
        RECT  17.300 1.420 17.530 3.780 ;
        RECT  17.110 1.420 17.300 1.650 ;
        RECT  16.655 2.795 17.300 3.025 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.440 1.945 9.955 2.175 ;
        RECT  8.425 1.945 8.440 2.595 ;
        RECT  8.195 1.945 8.425 2.635 ;
        RECT  8.135 2.365 8.195 2.635 ;
        RECT  6.390 2.365 8.135 2.595 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 2.050 15.505 2.280 ;
        RECT  12.170 1.845 12.400 2.280 ;
        RECT  12.095 1.845 12.170 2.075 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.090 -0.400 18.480 0.400 ;
        RECT  17.750 -0.400 18.090 0.960 ;
        RECT  16.810 -0.400 17.750 0.400 ;
        RECT  16.470 -0.400 16.810 0.960 ;
        RECT  15.465 -0.400 16.470 0.400 ;
        RECT  15.125 -0.400 15.465 0.950 ;
        RECT  14.185 -0.400 15.125 0.400 ;
        RECT  13.845 -0.400 14.185 0.950 ;
        RECT  12.905 -0.400 13.845 0.400 ;
        RECT  12.565 -0.400 12.905 0.895 ;
        RECT  4.680 -0.400 12.565 0.400 ;
        RECT  4.340 -0.400 4.680 0.575 ;
        RECT  3.120 -0.400 4.340 0.400 ;
        RECT  2.780 -0.400 3.120 0.575 ;
        RECT  1.800 -0.400 2.780 0.400 ;
        RECT  1.460 -0.400 1.800 0.960 ;
        RECT  0.520 -0.400 1.460 0.400 ;
        RECT  0.180 -0.400 0.520 0.950 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.745 4.640 18.480 5.440 ;
        RECT  17.295 4.465 17.745 5.440 ;
        RECT  16.335 4.640 17.295 5.440 ;
        RECT  15.995 4.090 16.335 5.440 ;
        RECT  15.030 4.640 15.995 5.440 ;
        RECT  14.690 4.090 15.030 5.440 ;
        RECT  13.750 4.640 14.690 5.440 ;
        RECT  13.410 4.090 13.750 5.440 ;
        RECT  12.425 4.640 13.410 5.440 ;
        RECT  12.085 4.465 12.425 5.440 ;
        RECT  10.865 4.640 12.085 5.440 ;
        RECT  10.525 4.465 10.865 5.440 ;
        RECT  4.480 4.640 10.525 5.440 ;
        RECT  4.140 4.465 4.480 5.440 ;
        RECT  3.120 4.640 4.140 5.440 ;
        RECT  2.780 4.465 3.120 5.440 ;
        RECT  1.800 4.640 2.780 5.440 ;
        RECT  1.460 4.090 1.800 5.440 ;
        RECT  0.520 4.640 1.460 5.440 ;
        RECT  0.180 4.090 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.160 2.095 16.755 2.325 ;
        RECT  15.930 2.095 16.160 2.765 ;
        RECT  13.490 1.490 16.105 1.720 ;
        RECT  11.640 2.535 15.930 2.765 ;
        RECT  12.300 3.005 15.675 3.235 ;
        RECT  13.205 1.360 13.490 1.720 ;
        RECT  12.230 1.360 13.205 1.590 ;
        RECT  12.070 3.005 12.300 3.680 ;
        RECT  12.000 0.715 12.230 1.590 ;
        RECT  10.705 3.450 12.070 3.680 ;
        RECT  11.110 0.715 12.000 0.945 ;
        RECT  11.570 2.535 11.640 3.125 ;
        RECT  11.340 1.390 11.570 3.125 ;
        RECT  11.285 2.895 11.340 3.125 ;
        RECT  10.880 0.715 11.110 1.645 ;
        RECT  10.705 1.415 10.880 1.645 ;
        RECT  10.475 1.415 10.705 4.215 ;
        RECT  8.445 1.415 10.475 1.645 ;
        RECT  8.020 3.985 10.475 4.215 ;
        RECT  7.790 3.680 8.020 4.215 ;
        RECT  5.385 3.680 7.790 3.910 ;
        RECT  5.160 0.665 7.425 0.895 ;
        RECT  4.940 4.145 7.040 4.375 ;
        RECT  5.155 3.535 5.385 3.910 ;
        RECT  4.930 0.665 5.160 1.040 ;
        RECT  2.905 3.535 5.155 3.765 ;
        RECT  3.745 1.515 4.975 1.745 ;
        RECT  4.710 4.005 4.940 4.375 ;
        RECT  2.875 0.810 4.930 1.040 ;
        RECT  2.440 4.005 4.710 4.235 ;
        RECT  3.515 1.515 3.745 3.080 ;
        RECT  2.680 2.180 2.905 3.765 ;
        RECT  2.645 0.810 2.875 1.645 ;
        RECT  2.675 2.070 2.680 3.765 ;
        RECT  0.930 2.070 2.675 2.410 ;
        RECT  0.695 1.415 2.645 1.645 ;
        RECT  2.210 2.795 2.440 4.235 ;
        RECT  0.695 2.795 2.210 3.025 ;
        RECT  0.465 1.415 0.695 3.025 ;
    END
END ADDHX4

MACRO ADDHX2
    CLASS CORE ;
    FOREIGN ADDHX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDHXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.715 1.285 5.945 1.645 ;
        RECT  4.240 2.830 5.860 3.170 ;
        RECT  3.515 1.340 5.715 1.570 ;
        RECT  3.745 2.885 4.240 3.170 ;
        RECT  3.265 2.885 3.745 3.195 ;
        RECT  3.320 1.285 3.515 1.570 ;
        RECT  3.265 1.285 3.320 1.625 ;
        RECT  3.035 1.285 3.265 3.195 ;
        RECT  2.980 1.285 3.035 1.625 ;
        RECT  3.015 2.810 3.035 3.195 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.080 1.360 11.505 1.700 ;
        RECT  11.005 1.360 11.080 1.845 ;
        RECT  11.015 2.630 11.070 3.080 ;
        RECT  11.005 2.630 11.015 3.195 ;
        RECT  10.775 1.470 11.005 3.195 ;
        RECT  10.730 2.630 10.775 3.080 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.145 1.840 5.485 2.180 ;
        RECT  5.065 1.840 5.145 2.125 ;
        RECT  4.835 1.845 5.065 2.125 ;
        RECT  4.100 1.895 4.835 2.125 ;
        RECT  3.870 1.895 4.100 2.600 ;
        RECT  3.760 2.260 3.870 2.600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.365 1.905 9.375 2.245 ;
        RECT  8.135 1.845 8.365 2.245 ;
        RECT  7.625 1.905 8.135 2.245 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.785 -0.400 11.880 0.400 ;
        RECT  10.445 -0.400 10.785 0.950 ;
        RECT  9.525 -0.400 10.445 0.400 ;
        RECT  9.185 -0.400 9.525 0.985 ;
        RECT  8.245 -0.400 9.185 0.400 ;
        RECT  7.905 -0.400 8.245 0.985 ;
        RECT  1.840 -0.400 7.905 0.400 ;
        RECT  1.500 -0.400 1.840 0.575 ;
        RECT  0.520 -0.400 1.500 0.400 ;
        RECT  0.180 -0.400 0.520 0.965 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.430 4.640 11.880 5.440 ;
        RECT  10.090 4.090 10.430 5.440 ;
        RECT  9.090 4.640 10.090 5.440 ;
        RECT  8.750 4.090 9.090 5.440 ;
        RECT  7.810 4.640 8.750 5.440 ;
        RECT  7.470 4.145 7.810 5.440 ;
        RECT  6.560 4.640 7.470 5.440 ;
        RECT  6.220 4.410 6.560 5.440 ;
        RECT  1.840 4.640 6.220 5.440 ;
        RECT  1.500 4.465 1.840 5.440 ;
        RECT  0.520 4.640 1.500 5.440 ;
        RECT  0.180 4.145 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.245 2.160 10.355 2.500 ;
        RECT  10.015 2.160 10.245 2.765 ;
        RECT  9.825 1.315 10.165 1.655 ;
        RECT  7.120 2.535 10.015 2.765 ;
        RECT  7.410 1.360 9.825 1.590 ;
        RECT  8.340 2.995 9.730 3.335 ;
        RECT  8.110 2.995 8.340 3.765 ;
        RECT  6.405 3.535 8.110 3.765 ;
        RECT  7.180 0.665 7.410 1.590 ;
        RECT  6.405 0.665 7.180 0.895 ;
        RECT  6.870 2.535 7.120 3.200 ;
        RECT  6.780 1.215 6.870 3.200 ;
        RECT  6.640 1.215 6.780 2.765 ;
        RECT  6.175 0.665 6.405 3.765 ;
        RECT  5.020 0.665 6.175 0.895 ;
        RECT  5.710 3.535 6.175 3.765 ;
        RECT  5.480 3.535 5.710 4.300 ;
        RECT  5.220 4.070 5.480 4.300 ;
        RECT  4.880 4.070 5.220 4.410 ;
        RECT  2.365 4.180 4.880 4.410 ;
        RECT  2.300 0.665 3.960 0.895 ;
        RECT  2.945 3.715 3.940 3.945 ;
        RECT  2.715 3.540 2.945 3.945 ;
        RECT  2.505 1.270 2.735 3.080 ;
        RECT  1.440 3.540 2.715 3.770 ;
        RECT  2.260 1.270 2.505 1.500 ;
        RECT  2.260 2.740 2.505 3.080 ;
        RECT  2.135 4.000 2.365 4.410 ;
        RECT  2.070 0.665 2.300 1.040 ;
        RECT  0.980 4.000 2.135 4.230 ;
        RECT  1.440 0.810 2.070 1.040 ;
        RECT  1.210 0.810 1.440 3.770 ;
        RECT  0.820 1.365 1.210 1.705 ;
        RECT  0.820 2.740 1.210 3.080 ;
        RECT  0.750 3.570 0.980 4.230 ;
        RECT  0.580 2.120 0.920 2.460 ;
        RECT  0.495 3.570 0.750 3.800 ;
        RECT  0.495 2.230 0.580 2.460 ;
        RECT  0.265 2.230 0.495 3.800 ;
    END
END ADDHX2

MACRO ADDHX1
    CLASS CORE ;
    FOREIGN ADDHX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDHXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.330 4.235 3.220 ;
        RECT  3.590 1.330 4.005 1.560 ;
        RECT  3.245 2.840 4.005 3.220 ;
        RECT  3.360 1.210 3.590 1.560 ;
        RECT  3.015 2.840 3.245 3.730 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.610 1.845 7.705 2.075 ;
        RECT  7.400 1.380 7.610 2.075 ;
        RECT  7.380 1.380 7.400 3.115 ;
        RECT  7.170 1.845 7.380 3.115 ;
        RECT  7.025 2.885 7.170 3.115 ;
        RECT  6.795 2.885 7.025 3.970 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 2.520 6.065 3.445 ;
        RECT  5.160 3.215 5.835 3.445 ;
        RECT  4.930 3.215 5.160 4.235 ;
        RECT  2.785 4.005 4.930 4.235 ;
        RECT  3.545 1.800 3.775 2.520 ;
        RECT  2.785 2.290 3.545 2.520 ;
        RECT  2.555 2.290 2.785 4.235 ;
        RECT  2.195 2.290 2.555 2.660 ;
        RECT  2.115 2.290 2.195 2.575 ;
        RECT  1.775 2.235 2.115 2.575 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.820 5.075 2.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.150 -0.400 7.920 0.400 ;
        RECT  6.920 -0.400 7.150 1.355 ;
        RECT  5.125 -0.400 6.920 0.400 ;
        RECT  6.815 1.125 6.920 1.355 ;
        RECT  6.585 1.125 6.815 1.720 ;
        RECT  4.785 -0.400 5.125 0.575 ;
        RECT  1.360 -0.400 4.785 0.400 ;
        RECT  1.020 -0.400 1.360 0.575 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.480 4.640 7.920 5.440 ;
        RECT  6.140 4.465 6.480 5.440 ;
        RECT  4.780 4.640 6.140 5.440 ;
        RECT  4.440 4.465 4.780 5.440 ;
        RECT  1.280 4.640 4.440 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.525 1.980 6.840 2.320 ;
        RECT  6.350 0.665 6.690 0.895 ;
        RECT  6.350 1.980 6.525 3.905 ;
        RECT  6.295 0.665 6.350 3.905 ;
        RECT  6.120 0.665 6.295 2.210 ;
        RECT  5.625 3.675 6.295 3.905 ;
        RECT  5.600 1.210 5.885 1.550 ;
        RECT  5.395 3.675 5.625 4.040 ;
        RECT  5.545 1.210 5.600 2.985 ;
        RECT  5.370 1.265 5.545 2.985 ;
        RECT  4.700 1.265 5.370 1.495 ;
        RECT  4.700 2.755 5.370 2.985 ;
        RECT  4.470 0.805 4.700 1.495 ;
        RECT  4.470 2.755 4.700 3.775 ;
        RECT  4.365 0.805 4.470 1.035 ;
        RECT  3.680 3.545 4.470 3.775 ;
        RECT  4.025 0.675 4.365 1.035 ;
        RECT  3.130 0.675 4.025 0.905 ;
        RECT  2.900 0.675 3.130 1.955 ;
        RECT  1.385 1.725 2.900 1.955 ;
        RECT  2.440 0.630 2.670 1.035 ;
        RECT  0.925 1.265 2.550 1.495 ;
        RECT  0.465 0.805 2.440 1.035 ;
        RECT  2.095 4.005 2.325 4.405 ;
        RECT  0.465 4.005 2.095 4.235 ;
        RECT  1.500 3.180 1.840 3.520 ;
        RECT  0.925 3.180 1.500 3.410 ;
        RECT  1.155 1.725 1.385 2.560 ;
        RECT  0.695 1.265 0.925 3.410 ;
        RECT  0.235 0.760 0.465 4.235 ;
    END
END ADDHX1

MACRO ADDFXL
    CLASS CORE ;
    FOREIGN ADDFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.570 1.285 13.645 1.515 ;
        RECT  13.460 1.285 13.570 1.845 ;
        RECT  13.460 2.635 13.570 3.605 ;
        RECT  13.230 1.285 13.460 3.605 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.005 2.380 12.325 2.660 ;
        RECT  11.985 1.430 12.005 2.660 ;
        RECT  11.755 1.430 11.985 3.135 ;
        RECT  11.665 1.430 11.755 1.770 ;
        RECT  11.645 2.795 11.755 3.135 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.220 1.820 9.485 2.050 ;
        RECT  8.990 1.820 9.220 3.220 ;
        RECT  8.600 2.865 8.990 3.220 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.040 0.760 2.380 ;
        RECT  0.420 2.040 0.445 2.635 ;
        RECT  0.215 2.150 0.420 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 2.350 4.835 2.690 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.770 -0.400 13.860 0.400 ;
        RECT  12.430 -0.400 12.770 1.615 ;
        RECT  10.080 -0.400 12.430 0.400 ;
        RECT  9.740 -0.400 10.080 0.575 ;
        RECT  4.725 -0.400 9.740 0.400 ;
        RECT  4.385 -0.400 4.725 0.900 ;
        RECT  1.285 -0.400 4.385 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.775 4.640 13.860 5.440 ;
        RECT  12.435 3.930 12.775 5.440 ;
        RECT  8.935 4.640 12.435 5.440 ;
        RECT  8.595 4.465 8.935 5.440 ;
        RECT  1.200 4.640 8.595 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.635 2.015 12.865 3.595 ;
        RECT  11.645 3.365 12.635 3.595 ;
        RECT  11.415 3.365 11.645 3.945 ;
        RECT  9.395 4.180 11.455 4.410 ;
        RECT  10.455 3.715 11.415 3.945 ;
        RECT  11.140 0.630 11.295 0.860 ;
        RECT  11.140 3.120 11.175 3.460 ;
        RECT  10.910 0.630 11.140 3.460 ;
        RECT  10.900 0.630 10.910 1.040 ;
        RECT  10.835 3.120 10.910 3.460 ;
        RECT  9.495 0.810 10.900 1.040 ;
        RECT  10.455 1.345 10.680 1.770 ;
        RECT  10.450 1.345 10.455 3.945 ;
        RECT  10.225 1.540 10.450 3.945 ;
        RECT  10.115 3.215 10.225 3.555 ;
        RECT  9.730 1.270 9.960 2.875 ;
        RECT  9.035 1.270 9.730 1.500 ;
        RECT  9.680 2.645 9.730 2.875 ;
        RECT  9.450 2.645 9.680 3.555 ;
        RECT  9.265 0.630 9.495 1.040 ;
        RECT  9.165 4.005 9.395 4.410 ;
        RECT  5.880 0.630 9.265 0.860 ;
        RECT  7.855 4.005 9.165 4.235 ;
        RECT  8.805 1.090 9.035 1.500 ;
        RECT  6.670 1.090 8.805 1.320 ;
        RECT  8.570 2.195 8.760 2.535 ;
        RECT  8.340 1.585 8.570 2.535 ;
        RECT  8.315 2.305 8.340 2.535 ;
        RECT  8.085 2.305 8.315 3.770 ;
        RECT  7.850 3.580 7.855 4.235 ;
        RECT  7.625 1.585 7.850 4.235 ;
        RECT  7.620 1.585 7.625 3.810 ;
        RECT  7.175 3.580 7.620 3.810 ;
        RECT  7.160 1.790 7.390 3.350 ;
        RECT  7.130 1.790 7.160 2.020 ;
        RECT  6.795 3.120 7.160 3.350 ;
        RECT  6.900 1.585 7.130 2.020 ;
        RECT  6.670 2.360 6.930 2.700 ;
        RECT  6.685 3.120 6.795 3.780 ;
        RECT  6.565 3.120 6.685 4.410 ;
        RECT  6.440 1.090 6.670 2.890 ;
        RECT  6.455 3.440 6.565 4.410 ;
        RECT  5.255 4.055 6.455 4.410 ;
        RECT  6.175 2.655 6.440 2.890 ;
        RECT  5.300 2.070 6.210 2.420 ;
        RECT  6.075 2.655 6.175 3.425 ;
        RECT  5.945 2.655 6.075 3.480 ;
        RECT  5.765 3.140 5.945 3.480 ;
        RECT  5.650 0.630 5.880 1.750 ;
        RECT  5.735 3.140 5.765 3.825 ;
        RECT  5.535 3.195 5.735 3.825 ;
        RECT  5.540 1.135 5.650 1.750 ;
        RECT  4.155 1.135 5.540 1.365 ;
        RECT  3.440 3.595 5.535 3.825 ;
        RECT  5.070 1.635 5.300 3.365 ;
        RECT  1.660 4.180 5.255 4.410 ;
        RECT  3.695 1.635 5.070 1.865 ;
        RECT  3.900 3.135 5.070 3.365 ;
        RECT  3.925 0.875 4.155 1.365 ;
        RECT  2.450 0.875 3.925 1.105 ;
        RECT  3.670 2.980 3.900 3.365 ;
        RECT  3.465 1.440 3.695 1.865 ;
        RECT  3.210 3.030 3.440 3.825 ;
        RECT  3.180 3.030 3.210 3.260 ;
        RECT  2.950 2.075 3.180 3.260 ;
        RECT  2.750 3.495 2.980 3.950 ;
        RECT  2.910 2.075 2.950 2.305 ;
        RECT  2.680 1.420 2.910 2.305 ;
        RECT  2.125 3.495 2.750 3.725 ;
        RECT  2.450 2.535 2.620 3.265 ;
        RECT  2.390 0.875 2.450 3.265 ;
        RECT  2.220 0.875 2.390 2.765 ;
        RECT  1.990 3.050 2.125 3.725 ;
        RECT  1.895 1.395 1.990 3.725 ;
        RECT  1.760 1.395 1.895 3.280 ;
        RECT  1.505 2.940 1.760 3.280 ;
        RECT  1.430 3.655 1.660 4.410 ;
        RECT  1.380 2.040 1.490 2.380 ;
        RECT  1.235 3.655 1.430 3.885 ;
        RECT  1.235 1.395 1.380 2.380 ;
        RECT  1.150 1.395 1.235 3.885 ;
        RECT  0.520 1.395 1.150 1.625 ;
        RECT  1.005 2.095 1.150 3.885 ;
        RECT  0.180 2.890 1.005 3.230 ;
        RECT  0.180 0.815 0.520 1.625 ;
    END
END ADDFXL

MACRO ADDFX4
    CLASS CORE ;
    FOREIGN ADDFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.720 1.395 13.935 3.155 ;
        RECT  13.595 1.395 13.720 3.220 ;
        RECT  13.340 1.820 13.595 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 1.395 12.655 3.155 ;
        RECT  12.315 1.395 12.400 3.220 ;
        RECT  12.020 1.820 12.315 3.220 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.220 1.820 9.485 2.050 ;
        RECT  8.990 1.820 9.220 3.220 ;
        RECT  8.600 2.865 8.990 3.220 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.040 0.760 2.380 ;
        RECT  0.420 2.040 0.445 2.635 ;
        RECT  0.215 2.150 0.420 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 2.350 4.835 2.690 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.575 -0.400 15.180 0.400 ;
        RECT  14.235 -0.400 14.575 1.005 ;
        RECT  13.295 -0.400 14.235 0.400 ;
        RECT  12.955 -0.400 13.295 1.005 ;
        RECT  12.015 -0.400 12.955 0.400 ;
        RECT  11.675 -0.400 12.015 1.005 ;
        RECT  10.080 -0.400 11.675 0.400 ;
        RECT  9.740 -0.400 10.080 0.575 ;
        RECT  4.725 -0.400 9.740 0.400 ;
        RECT  4.385 -0.400 4.725 0.905 ;
        RECT  1.285 -0.400 4.385 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.555 4.640 15.180 5.440 ;
        RECT  14.215 4.145 14.555 5.440 ;
        RECT  13.275 4.640 14.215 5.440 ;
        RECT  12.935 4.145 13.275 5.440 ;
        RECT  11.995 4.640 12.935 5.440 ;
        RECT  11.655 4.145 11.995 5.440 ;
        RECT  8.935 4.640 11.655 5.440 ;
        RECT  8.595 4.465 8.935 5.440 ;
        RECT  1.200 4.640 8.595 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.165 2.015 14.395 3.915 ;
        RECT  10.455 3.685 14.165 3.915 ;
        RECT  9.395 4.180 11.365 4.410 ;
        RECT  11.185 0.630 11.285 0.860 ;
        RECT  10.955 0.630 11.185 3.420 ;
        RECT  10.900 0.630 10.955 1.040 ;
        RECT  10.835 3.175 10.955 3.420 ;
        RECT  9.495 0.810 10.900 1.040 ;
        RECT  10.450 1.345 10.670 2.360 ;
        RECT  10.450 3.215 10.455 3.915 ;
        RECT  10.440 1.345 10.450 3.915 ;
        RECT  10.225 2.130 10.440 3.915 ;
        RECT  10.220 2.130 10.225 3.555 ;
        RECT  10.115 3.215 10.220 3.555 ;
        RECT  9.720 1.270 9.950 2.875 ;
        RECT  9.035 1.270 9.720 1.500 ;
        RECT  9.680 2.645 9.720 2.875 ;
        RECT  9.450 2.645 9.680 3.555 ;
        RECT  9.265 0.630 9.495 1.040 ;
        RECT  9.165 4.005 9.395 4.410 ;
        RECT  5.880 0.630 9.265 0.860 ;
        RECT  7.855 4.005 9.165 4.235 ;
        RECT  8.805 1.090 9.035 1.500 ;
        RECT  6.670 1.090 8.805 1.320 ;
        RECT  8.570 2.195 8.760 2.535 ;
        RECT  8.340 1.585 8.570 2.535 ;
        RECT  8.315 2.305 8.340 2.535 ;
        RECT  8.085 2.305 8.315 3.770 ;
        RECT  7.850 3.580 7.855 4.235 ;
        RECT  7.625 1.585 7.850 4.235 ;
        RECT  7.620 1.585 7.625 3.810 ;
        RECT  7.175 3.580 7.620 3.810 ;
        RECT  7.160 1.790 7.390 3.350 ;
        RECT  7.130 1.790 7.160 2.020 ;
        RECT  6.795 3.120 7.160 3.350 ;
        RECT  6.900 1.585 7.130 2.020 ;
        RECT  6.670 2.360 6.930 2.700 ;
        RECT  6.685 3.120 6.795 3.845 ;
        RECT  6.565 3.120 6.685 4.410 ;
        RECT  6.440 1.090 6.670 2.890 ;
        RECT  6.455 3.505 6.565 4.410 ;
        RECT  5.255 4.055 6.455 4.410 ;
        RECT  6.175 2.655 6.440 2.890 ;
        RECT  5.300 2.070 6.210 2.420 ;
        RECT  6.075 2.655 6.175 3.425 ;
        RECT  5.945 2.655 6.075 3.480 ;
        RECT  5.765 3.140 5.945 3.480 ;
        RECT  5.650 0.630 5.880 1.750 ;
        RECT  5.735 3.140 5.765 3.825 ;
        RECT  5.535 3.195 5.735 3.825 ;
        RECT  5.540 1.135 5.650 1.750 ;
        RECT  4.155 1.135 5.540 1.365 ;
        RECT  3.440 3.595 5.535 3.825 ;
        RECT  5.070 1.635 5.300 3.365 ;
        RECT  1.660 4.180 5.255 4.410 ;
        RECT  3.695 1.635 5.070 1.865 ;
        RECT  3.900 3.135 5.070 3.365 ;
        RECT  3.925 0.875 4.155 1.365 ;
        RECT  2.450 0.875 3.925 1.105 ;
        RECT  3.670 2.980 3.900 3.365 ;
        RECT  3.465 1.440 3.695 1.865 ;
        RECT  3.210 3.030 3.440 3.825 ;
        RECT  3.180 3.030 3.210 3.260 ;
        RECT  2.950 2.075 3.180 3.260 ;
        RECT  2.750 3.495 2.980 3.950 ;
        RECT  2.910 2.075 2.950 2.305 ;
        RECT  2.680 1.420 2.910 2.305 ;
        RECT  2.125 3.495 2.750 3.725 ;
        RECT  2.450 2.535 2.620 3.160 ;
        RECT  2.390 0.875 2.450 3.160 ;
        RECT  2.220 0.875 2.390 2.765 ;
        RECT  1.990 3.050 2.125 3.725 ;
        RECT  1.895 1.395 1.990 3.725 ;
        RECT  1.760 1.395 1.895 3.280 ;
        RECT  1.505 2.940 1.760 3.280 ;
        RECT  1.430 3.655 1.660 4.410 ;
        RECT  1.380 2.040 1.490 2.380 ;
        RECT  1.235 3.655 1.430 3.885 ;
        RECT  1.235 1.395 1.380 2.380 ;
        RECT  1.150 1.395 1.235 3.885 ;
        RECT  0.520 1.395 1.150 1.625 ;
        RECT  1.005 2.095 1.150 3.885 ;
        RECT  0.180 2.890 1.005 3.230 ;
        RECT  0.180 0.815 0.520 1.625 ;
    END
END ADDFX4

MACRO ADDFX2
    CLASS CORE ;
    FOREIGN ADDFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.325 1.285 13.370 1.780 ;
        RECT  13.325 2.795 13.355 3.135 ;
        RECT  13.095 1.285 13.325 3.135 ;
        RECT  13.030 1.285 13.095 1.780 ;
        RECT  13.015 2.795 13.095 3.135 ;
        RECT  12.755 1.285 13.030 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.760 1.430 12.005 1.770 ;
        RECT  11.760 2.795 11.985 3.135 ;
        RECT  11.530 1.430 11.760 3.135 ;
        RECT  11.435 2.405 11.530 2.635 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.220 1.820 9.485 2.050 ;
        RECT  8.990 1.820 9.220 3.220 ;
        RECT  8.600 2.865 8.990 3.220 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.040 0.760 2.380 ;
        RECT  0.420 2.040 0.445 2.635 ;
        RECT  0.215 2.150 0.420 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 2.350 4.835 2.690 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.690 -0.400 13.860 0.400 ;
        RECT  12.350 -0.400 12.690 0.575 ;
        RECT  10.080 -0.400 12.350 0.400 ;
        RECT  9.740 -0.400 10.080 0.575 ;
        RECT  4.725 -0.400 9.740 0.400 ;
        RECT  4.385 -0.400 4.725 0.900 ;
        RECT  1.285 -0.400 4.385 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.675 4.640 13.860 5.440 ;
        RECT  12.335 4.465 12.675 5.440 ;
        RECT  8.935 4.640 12.335 5.440 ;
        RECT  8.595 4.465 8.935 5.440 ;
        RECT  1.200 4.640 8.595 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.635 2.015 12.865 2.390 ;
        RECT  12.515 2.160 12.635 2.390 ;
        RECT  12.285 2.160 12.515 3.945 ;
        RECT  10.455 3.715 12.285 3.945 ;
        RECT  9.395 4.180 11.365 4.410 ;
        RECT  11.130 0.630 11.285 0.860 ;
        RECT  11.130 3.120 11.175 3.460 ;
        RECT  10.900 0.630 11.130 3.460 ;
        RECT  9.495 0.810 10.900 1.040 ;
        RECT  10.835 3.120 10.900 3.460 ;
        RECT  10.450 1.345 10.670 2.360 ;
        RECT  10.450 3.215 10.455 3.945 ;
        RECT  10.440 1.345 10.450 3.945 ;
        RECT  10.225 2.130 10.440 3.945 ;
        RECT  10.220 2.130 10.225 3.555 ;
        RECT  10.115 3.215 10.220 3.555 ;
        RECT  9.720 1.270 9.950 2.875 ;
        RECT  9.035 1.270 9.720 1.500 ;
        RECT  9.680 2.645 9.720 2.875 ;
        RECT  9.450 2.645 9.680 3.555 ;
        RECT  9.265 0.630 9.495 1.040 ;
        RECT  9.165 4.005 9.395 4.410 ;
        RECT  5.880 0.630 9.265 0.860 ;
        RECT  7.855 4.005 9.165 4.235 ;
        RECT  8.805 1.090 9.035 1.500 ;
        RECT  6.670 1.090 8.805 1.320 ;
        RECT  8.570 2.195 8.760 2.535 ;
        RECT  8.340 1.585 8.570 2.535 ;
        RECT  8.315 2.305 8.340 2.535 ;
        RECT  8.085 2.305 8.315 3.770 ;
        RECT  7.850 3.580 7.855 4.235 ;
        RECT  7.625 1.585 7.850 4.235 ;
        RECT  7.620 1.585 7.625 3.810 ;
        RECT  7.175 3.580 7.620 3.810 ;
        RECT  7.160 1.790 7.390 3.350 ;
        RECT  7.130 1.790 7.160 2.020 ;
        RECT  6.795 3.120 7.160 3.350 ;
        RECT  6.900 1.585 7.130 2.020 ;
        RECT  6.670 2.360 6.930 2.700 ;
        RECT  6.685 3.120 6.795 3.845 ;
        RECT  6.565 3.120 6.685 4.410 ;
        RECT  6.440 1.090 6.670 2.890 ;
        RECT  6.455 3.505 6.565 4.410 ;
        RECT  5.255 4.055 6.455 4.410 ;
        RECT  6.175 2.655 6.440 2.890 ;
        RECT  5.300 2.070 6.210 2.420 ;
        RECT  6.075 2.655 6.175 3.425 ;
        RECT  5.945 2.655 6.075 3.480 ;
        RECT  5.765 3.140 5.945 3.480 ;
        RECT  5.650 0.630 5.880 1.750 ;
        RECT  5.735 3.140 5.765 3.825 ;
        RECT  5.535 3.195 5.735 3.825 ;
        RECT  5.540 1.135 5.650 1.750 ;
        RECT  4.155 1.135 5.540 1.365 ;
        RECT  3.440 3.595 5.535 3.825 ;
        RECT  5.070 1.635 5.300 3.365 ;
        RECT  1.660 4.180 5.255 4.410 ;
        RECT  3.695 1.635 5.070 1.865 ;
        RECT  3.900 3.135 5.070 3.365 ;
        RECT  3.925 0.875 4.155 1.365 ;
        RECT  2.450 0.875 3.925 1.105 ;
        RECT  3.670 2.980 3.900 3.365 ;
        RECT  3.465 1.440 3.695 1.865 ;
        RECT  3.210 3.030 3.440 3.825 ;
        RECT  3.180 3.030 3.210 3.260 ;
        RECT  2.950 2.075 3.180 3.260 ;
        RECT  2.750 3.495 2.980 3.950 ;
        RECT  2.910 2.075 2.950 2.305 ;
        RECT  2.680 1.420 2.910 2.305 ;
        RECT  2.125 3.495 2.750 3.725 ;
        RECT  2.450 2.535 2.620 3.160 ;
        RECT  2.390 0.875 2.450 3.160 ;
        RECT  2.220 0.875 2.390 2.765 ;
        RECT  1.990 3.050 2.125 3.725 ;
        RECT  1.895 1.395 1.990 3.725 ;
        RECT  1.760 1.395 1.895 3.280 ;
        RECT  1.505 2.940 1.760 3.280 ;
        RECT  1.430 3.655 1.660 4.410 ;
        RECT  1.380 2.040 1.490 2.380 ;
        RECT  1.235 3.655 1.430 3.885 ;
        RECT  1.235 1.395 1.380 2.380 ;
        RECT  1.150 1.395 1.235 3.885 ;
        RECT  0.520 1.395 1.150 1.625 ;
        RECT  1.005 2.095 1.150 3.885 ;
        RECT  0.180 2.890 1.005 3.230 ;
        RECT  0.180 0.815 0.520 1.625 ;
    END
END ADDFX2

MACRO ADDFX1
    CLASS CORE ;
    FOREIGN ADDFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.570 1.285 13.645 1.515 ;
        RECT  13.460 1.285 13.570 1.845 ;
        RECT  13.460 2.635 13.570 3.605 ;
        RECT  13.230 1.285 13.460 3.605 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.005 2.380 12.325 2.660 ;
        RECT  11.985 1.430 12.005 2.660 ;
        RECT  11.755 1.430 11.985 3.135 ;
        RECT  11.665 1.430 11.755 1.770 ;
        RECT  11.645 2.795 11.755 3.135 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.220 1.820 9.485 2.050 ;
        RECT  8.990 1.820 9.220 3.220 ;
        RECT  8.600 2.865 8.990 3.220 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.040 0.760 2.380 ;
        RECT  0.420 2.040 0.445 2.635 ;
        RECT  0.215 2.150 0.420 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 2.350 4.835 2.690 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.770 -0.400 13.860 0.400 ;
        RECT  12.430 -0.400 12.770 1.615 ;
        RECT  10.080 -0.400 12.430 0.400 ;
        RECT  9.740 -0.400 10.080 0.575 ;
        RECT  4.725 -0.400 9.740 0.400 ;
        RECT  4.385 -0.400 4.725 0.900 ;
        RECT  1.285 -0.400 4.385 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.775 4.640 13.860 5.440 ;
        RECT  12.435 3.930 12.775 5.440 ;
        RECT  8.935 4.640 12.435 5.440 ;
        RECT  8.595 4.465 8.935 5.440 ;
        RECT  1.200 4.640 8.595 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.635 2.015 12.865 3.595 ;
        RECT  11.645 3.365 12.635 3.595 ;
        RECT  11.415 3.365 11.645 3.945 ;
        RECT  9.395 4.180 11.455 4.410 ;
        RECT  10.455 3.715 11.415 3.945 ;
        RECT  11.140 0.630 11.295 0.860 ;
        RECT  11.140 3.120 11.175 3.460 ;
        RECT  10.910 0.630 11.140 3.460 ;
        RECT  10.900 0.630 10.910 1.040 ;
        RECT  10.835 3.120 10.910 3.460 ;
        RECT  9.495 0.810 10.900 1.040 ;
        RECT  10.455 1.345 10.680 1.770 ;
        RECT  10.450 1.345 10.455 3.945 ;
        RECT  10.225 1.540 10.450 3.945 ;
        RECT  10.115 3.215 10.225 3.555 ;
        RECT  9.730 1.270 9.960 2.875 ;
        RECT  9.035 1.270 9.730 1.500 ;
        RECT  9.680 2.645 9.730 2.875 ;
        RECT  9.450 2.645 9.680 3.555 ;
        RECT  9.265 0.630 9.495 1.040 ;
        RECT  9.165 4.005 9.395 4.410 ;
        RECT  5.880 0.630 9.265 0.860 ;
        RECT  7.855 4.005 9.165 4.235 ;
        RECT  8.805 1.090 9.035 1.500 ;
        RECT  6.670 1.090 8.805 1.320 ;
        RECT  8.570 2.195 8.760 2.535 ;
        RECT  8.340 1.585 8.570 2.535 ;
        RECT  8.315 2.305 8.340 2.535 ;
        RECT  8.085 2.305 8.315 3.770 ;
        RECT  7.850 3.580 7.855 4.235 ;
        RECT  7.625 1.585 7.850 4.235 ;
        RECT  7.620 1.585 7.625 3.810 ;
        RECT  7.175 3.580 7.620 3.810 ;
        RECT  7.160 1.790 7.390 3.350 ;
        RECT  7.130 1.790 7.160 2.020 ;
        RECT  6.795 3.120 7.160 3.350 ;
        RECT  6.900 1.585 7.130 2.020 ;
        RECT  6.670 2.360 6.930 2.700 ;
        RECT  6.685 3.120 6.795 3.780 ;
        RECT  6.565 3.120 6.685 4.410 ;
        RECT  6.440 1.090 6.670 2.890 ;
        RECT  6.455 3.440 6.565 4.410 ;
        RECT  5.255 4.055 6.455 4.410 ;
        RECT  6.175 2.655 6.440 2.890 ;
        RECT  5.300 2.070 6.210 2.420 ;
        RECT  6.075 2.655 6.175 3.425 ;
        RECT  5.945 2.655 6.075 3.480 ;
        RECT  5.765 3.140 5.945 3.480 ;
        RECT  5.650 0.630 5.880 1.750 ;
        RECT  5.735 3.140 5.765 3.825 ;
        RECT  5.535 3.195 5.735 3.825 ;
        RECT  5.540 1.135 5.650 1.750 ;
        RECT  4.155 1.135 5.540 1.365 ;
        RECT  3.440 3.595 5.535 3.825 ;
        RECT  5.070 1.635 5.300 3.365 ;
        RECT  1.660 4.180 5.255 4.410 ;
        RECT  3.695 1.635 5.070 1.865 ;
        RECT  3.900 3.135 5.070 3.365 ;
        RECT  3.925 0.875 4.155 1.365 ;
        RECT  2.450 0.875 3.925 1.105 ;
        RECT  3.670 2.980 3.900 3.365 ;
        RECT  3.465 1.440 3.695 1.865 ;
        RECT  3.210 3.030 3.440 3.825 ;
        RECT  3.180 3.030 3.210 3.260 ;
        RECT  2.950 2.075 3.180 3.260 ;
        RECT  2.750 3.495 2.980 3.950 ;
        RECT  2.910 2.075 2.950 2.305 ;
        RECT  2.680 1.420 2.910 2.305 ;
        RECT  2.125 3.495 2.750 3.725 ;
        RECT  2.450 2.535 2.620 3.265 ;
        RECT  2.390 0.875 2.450 3.265 ;
        RECT  2.220 0.875 2.390 2.765 ;
        RECT  1.990 3.050 2.125 3.725 ;
        RECT  1.895 1.395 1.990 3.725 ;
        RECT  1.760 1.395 1.895 3.280 ;
        RECT  1.505 2.940 1.760 3.280 ;
        RECT  1.430 3.655 1.660 4.410 ;
        RECT  1.380 2.040 1.490 2.380 ;
        RECT  1.235 3.655 1.430 3.885 ;
        RECT  1.235 1.395 1.380 2.380 ;
        RECT  1.150 1.395 1.235 3.885 ;
        RECT  0.520 1.395 1.150 1.625 ;
        RECT  1.005 2.095 1.150 3.885 ;
        RECT  0.180 2.890 1.005 3.230 ;
        RECT  0.180 0.815 0.520 1.625 ;
    END
END ADDFX1

MACRO ADDFHXL
    CLASS CORE ;
    FOREIGN ADDFHXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.230 1.285 14.340 2.100 ;
        RECT  14.230 3.080 14.340 3.420 ;
        RECT  14.000 1.285 14.230 3.420 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.725 1.285 12.865 1.625 ;
        RECT  12.725 3.080 12.780 3.420 ;
        RECT  12.495 1.285 12.725 3.420 ;
        RECT  12.440 2.940 12.495 3.420 ;
        RECT  12.090 2.940 12.440 3.220 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.360 2.675 11.745 3.220 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 2.805 6.540 3.145 ;
        RECT  6.385 2.660 6.490 3.145 ;
        RECT  6.155 2.405 6.385 3.145 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 2.085 1.180 2.670 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.625 -0.400 14.520 0.400 ;
        RECT  13.285 -0.400 13.625 0.575 ;
        RECT  12.255 -0.400 13.285 0.400 ;
        RECT  11.915 -0.400 12.255 0.575 ;
        RECT  6.955 -0.400 11.915 0.400 ;
        RECT  6.615 -0.400 6.955 0.575 ;
        RECT  1.320 -0.400 6.615 0.400 ;
        RECT  0.980 -0.400 1.320 0.575 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.560 4.640 14.520 5.440 ;
        RECT  13.220 4.465 13.560 5.440 ;
        RECT  10.940 4.640 13.220 5.440 ;
        RECT  10.600 4.465 10.940 5.440 ;
        RECT  6.160 4.640 10.600 5.440 ;
        RECT  5.820 4.465 6.160 5.440 ;
        RECT  1.240 4.640 5.820 5.440 ;
        RECT  0.900 3.760 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.420 2.400 13.760 2.740 ;
        RECT  13.240 2.510 13.420 2.740 ;
        RECT  13.010 2.510 13.240 4.230 ;
        RECT  11.680 0.810 13.085 1.040 ;
        RECT  9.660 4.000 13.010 4.230 ;
        RECT  11.820 1.355 12.160 1.695 ;
        RECT  10.920 3.450 11.915 3.680 ;
        RECT  11.220 1.465 11.820 1.695 ;
        RECT  11.450 0.630 11.680 1.040 ;
        RECT  8.940 0.630 11.450 0.860 ;
        RECT  10.990 1.090 11.220 2.425 ;
        RECT  9.400 1.090 10.990 1.320 ;
        RECT  10.920 2.195 10.990 2.425 ;
        RECT  10.690 2.195 10.920 3.680 ;
        RECT  10.460 1.550 10.760 1.780 ;
        RECT  10.230 1.550 10.460 3.675 ;
        RECT  10.040 3.335 10.230 3.675 ;
        RECT  9.860 1.550 9.995 1.780 ;
        RECT  9.660 1.550 9.860 2.760 ;
        RECT  9.630 1.550 9.660 4.230 ;
        RECT  9.430 2.530 9.630 4.230 ;
        RECT  9.320 3.545 9.430 3.885 ;
        RECT  9.170 1.090 9.400 1.780 ;
        RECT  8.885 1.550 9.170 1.780 ;
        RECT  8.710 0.630 8.940 1.320 ;
        RECT  8.655 1.550 8.885 3.885 ;
        RECT  8.420 1.090 8.710 1.320 ;
        RECT  7.960 0.630 8.475 0.860 ;
        RECT  8.190 1.090 8.420 3.830 ;
        RECT  8.120 3.600 8.190 3.830 ;
        RECT  7.780 3.600 8.120 3.940 ;
        RECT  7.730 0.630 7.960 3.130 ;
        RECT  6.385 0.805 7.730 1.035 ;
        RECT  7.640 2.755 7.730 3.130 ;
        RECT  7.410 1.265 7.500 1.605 ;
        RECT  7.180 1.265 7.410 3.620 ;
        RECT  5.815 3.390 7.180 3.620 ;
        RECT  6.720 1.325 6.950 2.340 ;
        RECT  5.920 1.325 6.720 1.555 ;
        RECT  6.155 0.630 6.385 1.035 ;
        RECT  4.430 0.630 6.155 0.860 ;
        RECT  5.690 1.090 5.920 1.555 ;
        RECT  5.585 2.175 5.815 3.620 ;
        RECT  4.890 1.090 5.690 1.320 ;
        RECT  5.350 1.600 5.460 1.940 ;
        RECT  5.120 1.600 5.350 4.410 ;
        RECT  2.190 4.180 5.120 4.410 ;
        RECT  4.810 1.090 4.890 1.885 ;
        RECT  4.660 1.090 4.810 3.950 ;
        RECT  4.580 1.655 4.660 3.950 ;
        RECT  2.965 3.720 4.580 3.950 ;
        RECT  4.350 0.630 4.430 1.420 ;
        RECT  4.200 0.630 4.350 3.465 ;
        RECT  4.120 1.040 4.200 3.465 ;
        RECT  3.710 1.090 3.765 1.430 ;
        RECT  3.630 0.630 3.710 1.430 ;
        RECT  3.630 3.125 3.685 3.465 ;
        RECT  3.400 0.630 3.630 3.465 ;
        RECT  1.810 0.630 3.400 0.860 ;
        RECT  3.345 3.125 3.400 3.465 ;
        RECT  2.910 1.090 3.045 1.430 ;
        RECT  2.910 3.180 2.965 3.950 ;
        RECT  2.735 1.090 2.910 3.950 ;
        RECT  2.680 1.090 2.735 3.520 ;
        RECT  2.625 3.180 2.680 3.520 ;
        RECT  2.190 1.090 2.270 3.475 ;
        RECT  2.040 1.090 2.190 4.410 ;
        RECT  1.960 3.100 2.040 4.410 ;
        RECT  1.580 0.630 1.810 1.035 ;
        RECT  1.715 2.345 1.780 2.715 ;
        RECT  1.485 1.555 1.715 3.165 ;
        RECT  0.520 0.805 1.580 1.035 ;
        RECT  0.870 1.555 1.485 1.785 ;
        RECT  0.870 2.935 1.485 3.165 ;
        RECT  0.640 1.310 0.870 1.785 ;
        RECT  0.640 2.935 0.870 3.300 ;
        RECT  0.410 0.665 0.520 1.035 ;
        RECT  0.410 3.760 0.520 4.100 ;
        RECT  0.180 0.665 0.410 4.100 ;
    END
END ADDFHXL

MACRO ADDFHX4
    CLASS CORE ;
    FOREIGN ADDFHX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFHXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.150 1.820 22.300 3.220 ;
        RECT  21.920 1.400 22.150 3.220 ;
        RECT  21.710 1.400 21.920 1.740 ;
        RECT  21.710 2.820 21.920 3.160 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.830 1.820 20.980 3.220 ;
        RECT  20.600 1.455 20.830 3.220 ;
        RECT  20.430 1.455 20.600 1.685 ;
        RECT  20.425 2.820 20.600 3.160 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.995 2.380 19.660 2.765 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 2.665 14.070 3.005 ;
        RECT  13.415 2.665 13.645 3.195 ;
        RECT  12.790 2.665 13.415 3.005 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 1.820 1.245 2.400 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.690 -0.400 23.100 0.400 ;
        RECT  22.350 -0.400 22.690 1.040 ;
        RECT  21.410 -0.400 22.350 0.400 ;
        RECT  21.070 -0.400 21.410 1.040 ;
        RECT  20.050 -0.400 21.070 0.400 ;
        RECT  19.710 -0.400 20.050 0.575 ;
        RECT  13.580 -0.400 19.710 0.400 ;
        RECT  13.240 -0.400 13.580 0.575 ;
        RECT  3.270 -0.400 13.240 0.400 ;
        RECT  2.930 -0.400 3.270 0.575 ;
        RECT  1.250 -0.400 2.930 0.400 ;
        RECT  0.910 -0.400 1.250 0.575 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.695 4.640 23.100 5.440 ;
        RECT  22.355 4.085 22.695 5.440 ;
        RECT  21.410 4.640 22.355 5.440 ;
        RECT  21.070 4.085 21.410 5.440 ;
        RECT  20.125 4.640 21.070 5.440 ;
        RECT  19.785 4.090 20.125 5.440 ;
        RECT  18.815 4.640 19.785 5.440 ;
        RECT  18.365 4.465 18.815 5.440 ;
        RECT  14.090 4.640 18.365 5.440 ;
        RECT  13.750 4.010 14.090 5.440 ;
        RECT  12.650 4.640 13.750 5.440 ;
        RECT  12.310 4.010 12.650 5.440 ;
        RECT  3.660 4.640 12.310 5.440 ;
        RECT  3.320 3.765 3.660 5.440 ;
        RECT  1.445 4.640 3.320 5.440 ;
        RECT  1.105 4.000 1.445 5.440 ;
        RECT  0.000 4.640 1.105 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.440 2.210 21.625 2.580 ;
        RECT  21.210 2.210 21.440 3.835 ;
        RECT  17.265 3.605 21.210 3.835 ;
        RECT  20.305 2.025 20.360 2.365 ;
        RECT  20.020 1.915 20.305 2.365 ;
        RECT  19.910 1.915 20.020 2.145 ;
        RECT  19.680 1.005 19.910 2.145 ;
        RECT  19.055 1.005 19.680 1.235 ;
        RECT  18.590 1.495 19.450 1.725 ;
        RECT  18.590 3.045 19.365 3.275 ;
        RECT  18.825 0.630 19.055 1.235 ;
        RECT  15.965 0.630 18.825 0.860 ;
        RECT  18.360 1.090 18.590 3.275 ;
        RECT  16.490 1.090 18.360 1.320 ;
        RECT  18.165 2.305 18.360 2.670 ;
        RECT  17.930 1.550 18.130 1.780 ;
        RECT  17.930 2.990 17.985 3.330 ;
        RECT  17.700 1.550 17.930 3.330 ;
        RECT  17.645 2.990 17.700 3.330 ;
        RECT  17.210 1.550 17.405 1.780 ;
        RECT  17.210 3.295 17.265 4.105 ;
        RECT  16.980 1.550 17.210 4.105 ;
        RECT  16.925 3.295 16.980 4.105 ;
        RECT  16.490 3.155 16.545 3.965 ;
        RECT  16.260 1.090 16.490 3.965 ;
        RECT  16.205 3.155 16.260 3.965 ;
        RECT  15.910 0.630 15.965 1.520 ;
        RECT  15.680 0.630 15.910 3.430 ;
        RECT  15.625 0.700 15.680 1.520 ;
        RECT  15.660 3.200 15.680 3.430 ;
        RECT  15.320 3.200 15.660 4.020 ;
        RECT  15.165 0.635 15.395 2.880 ;
        RECT  15.150 0.635 15.165 1.035 ;
        RECT  12.745 0.805 15.150 1.035 ;
        RECT  14.810 1.460 14.935 3.680 ;
        RECT  14.705 1.460 14.810 4.310 ;
        RECT  14.340 1.460 14.705 1.690 ;
        RECT  14.470 3.450 14.705 4.310 ;
        RECT  14.245 1.920 14.475 2.290 ;
        RECT  13.370 3.450 14.470 3.680 ;
        RECT  14.000 1.350 14.340 1.690 ;
        RECT  13.260 1.920 14.245 2.150 ;
        RECT  13.030 3.450 13.370 4.310 ;
        RECT  13.030 1.265 13.260 2.150 ;
        RECT  12.195 1.265 13.030 1.495 ;
        RECT  12.195 3.450 13.030 3.680 ;
        RECT  12.195 1.725 12.780 1.955 ;
        RECT  12.515 0.660 12.745 1.035 ;
        RECT  9.705 0.660 12.515 0.890 ;
        RECT  11.965 1.130 12.195 1.495 ;
        RECT  11.965 1.725 12.195 3.780 ;
        RECT  10.165 1.130 11.965 1.360 ;
        RECT  11.505 1.595 11.735 4.295 ;
        RECT  10.395 1.595 11.505 1.825 ;
        RECT  9.970 4.065 11.505 4.295 ;
        RECT  11.035 2.060 11.265 3.815 ;
        RECT  10.165 2.060 11.035 2.290 ;
        RECT  7.240 3.585 11.035 3.815 ;
        RECT  10.580 3.100 10.785 3.330 ;
        RECT  10.350 2.525 10.580 3.330 ;
        RECT  9.705 2.525 10.350 2.755 ;
        RECT  9.935 1.130 10.165 2.290 ;
        RECT  9.685 4.065 9.970 4.340 ;
        RECT  9.475 0.630 9.705 2.755 ;
        RECT  4.380 4.110 9.685 4.340 ;
        RECT  9.190 3.095 9.480 3.325 ;
        RECT  8.340 0.630 9.475 0.860 ;
        RECT  8.960 1.260 9.190 3.325 ;
        RECT  8.720 1.260 8.960 1.490 ;
        RECT  7.815 3.095 8.960 3.325 ;
        RECT  8.285 2.635 8.720 2.865 ;
        RECT  8.285 0.630 8.340 1.330 ;
        RECT  8.110 0.630 8.285 2.865 ;
        RECT  8.055 0.990 8.110 2.865 ;
        RECT  8.000 0.990 8.055 1.330 ;
        RECT  7.585 1.950 7.815 3.325 ;
        RECT  7.565 0.990 7.620 1.330 ;
        RECT  7.565 1.950 7.585 2.180 ;
        RECT  7.510 0.990 7.565 2.180 ;
        RECT  7.335 0.630 7.510 2.180 ;
        RECT  7.280 0.630 7.335 1.330 ;
        RECT  6.175 0.630 7.280 0.860 ;
        RECT  7.185 3.045 7.240 3.865 ;
        RECT  6.980 2.460 7.185 3.865 ;
        RECT  6.955 1.185 6.980 3.865 ;
        RECT  6.750 1.185 6.955 2.690 ;
        RECT  6.900 3.045 6.955 3.865 ;
        RECT  5.045 3.635 6.900 3.865 ;
        RECT  6.560 1.185 6.750 1.415 ;
        RECT  6.390 3.095 6.520 3.325 ;
        RECT  6.160 2.400 6.390 3.325 ;
        RECT  6.120 0.630 6.175 1.130 ;
        RECT  6.120 2.400 6.160 2.630 ;
        RECT  5.890 0.630 6.120 2.630 ;
        RECT  5.835 0.630 5.890 1.130 ;
        RECT  3.735 0.630 5.835 0.860 ;
        RECT  5.510 3.100 5.820 3.330 ;
        RECT  5.480 1.605 5.510 3.330 ;
        RECT  5.425 1.550 5.480 3.330 ;
        RECT  5.280 1.090 5.425 3.330 ;
        RECT  5.195 1.090 5.280 1.920 ;
        RECT  4.200 1.090 5.195 1.320 ;
        RECT  5.140 1.550 5.195 1.890 ;
        RECT  4.815 2.505 5.045 3.865 ;
        RECT  4.695 2.505 4.815 2.735 ;
        RECT  4.465 1.550 4.695 2.735 ;
        RECT  4.150 3.100 4.380 4.340 ;
        RECT  4.030 1.090 4.200 1.685 ;
        RECT  4.040 3.100 4.150 3.985 ;
        RECT  3.780 3.100 4.040 3.530 ;
        RECT  3.970 1.090 4.030 1.740 ;
        RECT  3.780 1.400 3.970 1.740 ;
        RECT  3.690 1.400 3.780 3.530 ;
        RECT  3.505 0.630 3.735 1.040 ;
        RECT  3.550 1.455 3.690 3.530 ;
        RECT  2.710 1.455 3.550 1.685 ;
        RECT  2.940 3.300 3.550 3.530 ;
        RECT  0.520 0.810 3.505 1.040 ;
        RECT  2.850 2.090 3.190 2.430 ;
        RECT  2.600 3.300 2.940 3.640 ;
        RECT  1.955 2.145 2.850 2.375 ;
        RECT  2.370 1.400 2.710 1.740 ;
        RECT  1.965 4.055 2.400 4.285 ;
        RECT  1.955 1.460 2.010 1.800 ;
        RECT  1.735 3.450 1.965 4.285 ;
        RECT  1.785 1.460 1.955 2.375 ;
        RECT  1.785 2.740 1.840 3.080 ;
        RECT  1.725 1.460 1.785 3.080 ;
        RECT  0.520 3.450 1.735 3.680 ;
        RECT  1.670 1.460 1.725 1.800 ;
        RECT  1.555 2.145 1.725 3.080 ;
        RECT  1.500 2.740 1.555 3.080 ;
        RECT  0.465 0.810 0.520 1.630 ;
        RECT  0.465 2.830 0.520 4.250 ;
        RECT  0.290 0.810 0.465 4.250 ;
        RECT  0.235 1.290 0.290 4.250 ;
        RECT  0.180 1.290 0.235 1.630 ;
        RECT  0.180 2.830 0.235 4.250 ;
    END
END ADDFHX4

MACRO ADDFHX2
    CLASS CORE ;
    FOREIGN ADDFHX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFHXL ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.050 0.920 22.230 2.075 ;
        RECT  22.050 2.635 22.105 4.025 ;
        RECT  21.890 0.920 22.050 4.025 ;
        RECT  21.820 1.500 21.890 4.025 ;
        RECT  21.765 2.745 21.820 4.025 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.790 1.390 20.970 1.730 ;
        RECT  20.630 1.390 20.790 3.195 ;
        RECT  20.560 1.445 20.630 3.195 ;
        RECT  20.015 2.965 20.560 3.195 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.995 2.295 19.660 2.725 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 2.665 14.070 3.005 ;
        RECT  13.415 2.665 13.645 3.195 ;
        RECT  12.790 2.665 13.415 3.005 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 1.820 1.245 2.400 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.510 -0.400 22.440 0.400 ;
        RECT  21.170 -0.400 21.510 0.950 ;
        RECT  20.210 -0.400 21.170 0.400 ;
        RECT  19.870 -0.400 20.210 0.575 ;
        RECT  13.580 -0.400 19.870 0.400 ;
        RECT  13.240 -0.400 13.580 0.575 ;
        RECT  3.350 -0.400 13.240 0.400 ;
        RECT  3.010 -0.400 3.350 0.575 ;
        RECT  1.330 -0.400 3.010 0.400 ;
        RECT  0.990 -0.400 1.330 0.575 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.385 4.640 22.440 5.440 ;
        RECT  21.045 4.085 21.385 5.440 ;
        RECT  20.125 4.640 21.045 5.440 ;
        RECT  19.785 4.085 20.125 5.440 ;
        RECT  18.790 4.640 19.785 5.440 ;
        RECT  18.385 4.465 18.790 5.440 ;
        RECT  14.090 4.640 18.385 5.440 ;
        RECT  13.750 4.010 14.090 5.440 ;
        RECT  12.650 4.640 13.750 5.440 ;
        RECT  12.310 4.010 12.650 5.440 ;
        RECT  3.660 4.640 12.310 5.440 ;
        RECT  3.320 3.765 3.660 5.440 ;
        RECT  1.445 4.640 3.320 5.440 ;
        RECT  1.105 4.000 1.445 5.440 ;
        RECT  0.000 4.640 1.105 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.020 2.210 21.250 3.835 ;
        RECT  17.265 3.605 21.020 3.835 ;
        RECT  20.075 1.005 20.305 2.430 ;
        RECT  19.055 1.005 20.075 1.235 ;
        RECT  18.590 1.495 19.450 1.725 ;
        RECT  18.590 3.125 19.365 3.355 ;
        RECT  18.825 0.630 19.055 1.235 ;
        RECT  15.910 0.630 18.825 0.860 ;
        RECT  18.360 1.090 18.590 3.355 ;
        RECT  16.490 1.090 18.360 1.320 ;
        RECT  18.165 2.305 18.360 2.670 ;
        RECT  17.930 1.550 18.130 1.780 ;
        RECT  17.930 3.030 17.985 3.370 ;
        RECT  17.700 1.550 17.930 3.370 ;
        RECT  17.645 3.030 17.700 3.370 ;
        RECT  17.210 1.550 17.405 1.780 ;
        RECT  17.210 3.295 17.265 4.105 ;
        RECT  16.980 1.550 17.210 4.105 ;
        RECT  16.925 3.295 16.980 4.105 ;
        RECT  16.490 3.155 16.545 3.965 ;
        RECT  16.260 1.090 16.490 3.965 ;
        RECT  16.205 3.155 16.260 3.965 ;
        RECT  15.680 0.630 15.910 3.350 ;
        RECT  15.660 3.120 15.680 3.350 ;
        RECT  15.375 3.120 15.660 4.095 ;
        RECT  15.165 0.635 15.395 2.880 ;
        RECT  15.320 3.275 15.375 4.095 ;
        RECT  15.150 0.635 15.165 1.035 ;
        RECT  12.745 0.805 15.150 1.035 ;
        RECT  14.755 1.405 14.935 3.050 ;
        RECT  14.755 3.440 14.810 4.260 ;
        RECT  14.705 1.405 14.755 4.260 ;
        RECT  14.340 1.405 14.705 1.635 ;
        RECT  14.525 2.820 14.705 4.260 ;
        RECT  14.470 3.440 14.525 4.260 ;
        RECT  14.245 1.920 14.475 2.290 ;
        RECT  13.370 3.460 14.470 3.690 ;
        RECT  14.000 1.350 14.340 1.690 ;
        RECT  13.260 1.920 14.245 2.150 ;
        RECT  13.030 3.460 13.370 4.305 ;
        RECT  13.030 1.265 13.260 2.150 ;
        RECT  12.195 1.265 13.030 1.495 ;
        RECT  12.195 3.460 13.030 3.690 ;
        RECT  12.195 1.725 12.780 1.955 ;
        RECT  12.515 0.660 12.745 1.035 ;
        RECT  9.705 0.660 12.515 0.890 ;
        RECT  11.965 1.130 12.195 1.495 ;
        RECT  11.965 1.725 12.195 3.780 ;
        RECT  10.165 1.130 11.965 1.360 ;
        RECT  11.505 1.595 11.735 4.295 ;
        RECT  10.395 1.595 11.505 1.825 ;
        RECT  9.970 4.065 11.505 4.295 ;
        RECT  11.035 2.060 11.265 3.820 ;
        RECT  10.165 2.060 11.035 2.290 ;
        RECT  7.185 3.590 11.035 3.820 ;
        RECT  10.580 3.100 10.785 3.330 ;
        RECT  10.350 2.525 10.580 3.330 ;
        RECT  9.705 2.525 10.350 2.755 ;
        RECT  9.935 1.130 10.165 2.290 ;
        RECT  9.685 4.065 9.970 4.410 ;
        RECT  9.475 0.630 9.705 2.755 ;
        RECT  4.395 4.180 9.685 4.410 ;
        RECT  9.190 3.095 9.480 3.325 ;
        RECT  8.285 0.630 9.475 0.860 ;
        RECT  8.960 1.260 9.190 3.325 ;
        RECT  8.720 1.260 8.960 1.490 ;
        RECT  7.650 3.095 8.960 3.325 ;
        RECT  8.285 2.635 8.720 2.865 ;
        RECT  8.055 0.630 8.285 2.865 ;
        RECT  7.565 1.230 7.650 3.325 ;
        RECT  7.420 0.630 7.565 3.325 ;
        RECT  7.335 0.630 7.420 1.460 ;
        RECT  6.120 0.630 7.335 0.860 ;
        RECT  6.955 1.875 7.185 3.860 ;
        RECT  6.845 1.875 6.955 2.105 ;
        RECT  5.045 3.630 6.955 3.860 ;
        RECT  6.615 1.130 6.845 2.105 ;
        RECT  6.410 3.040 6.520 3.380 ;
        RECT  6.180 2.400 6.410 3.380 ;
        RECT  6.120 2.400 6.180 2.630 ;
        RECT  5.890 0.630 6.120 2.630 ;
        RECT  3.815 0.630 5.890 0.860 ;
        RECT  5.590 3.045 5.820 3.385 ;
        RECT  5.480 1.090 5.590 3.385 ;
        RECT  5.360 1.090 5.480 3.330 ;
        RECT  4.280 1.090 5.360 1.320 ;
        RECT  5.275 1.550 5.360 1.920 ;
        RECT  4.815 2.505 5.045 3.860 ;
        RECT  4.775 2.505 4.815 2.735 ;
        RECT  4.545 1.550 4.775 2.735 ;
        RECT  4.165 3.295 4.395 4.410 ;
        RECT  4.050 1.090 4.280 1.555 ;
        RECT  4.025 3.295 4.165 3.580 ;
        RECT  3.780 1.325 4.050 1.555 ;
        RECT  3.780 3.295 4.025 3.525 ;
        RECT  3.585 0.630 3.815 1.040 ;
        RECT  3.550 1.325 3.780 3.525 ;
        RECT  0.520 0.810 3.585 1.040 ;
        RECT  2.790 1.325 3.550 1.555 ;
        RECT  2.950 3.295 3.550 3.525 ;
        RECT  2.930 2.090 3.270 2.430 ;
        RECT  2.580 3.295 2.950 3.580 ;
        RECT  2.035 2.145 2.930 2.375 ;
        RECT  2.450 1.270 2.790 1.610 ;
        RECT  1.965 4.055 2.400 4.285 ;
        RECT  2.035 1.460 2.090 1.800 ;
        RECT  1.840 1.460 2.035 2.375 ;
        RECT  1.735 3.450 1.965 4.285 ;
        RECT  1.805 1.460 1.840 3.080 ;
        RECT  1.750 1.460 1.805 1.800 ;
        RECT  1.610 2.145 1.805 3.080 ;
        RECT  0.520 3.450 1.735 3.680 ;
        RECT  1.500 2.740 1.610 3.080 ;
        RECT  0.465 0.810 0.520 1.550 ;
        RECT  0.465 2.830 0.520 4.250 ;
        RECT  0.290 0.810 0.465 4.250 ;
        RECT  0.235 1.210 0.290 4.250 ;
        RECT  0.180 1.210 0.235 1.550 ;
        RECT  0.180 2.830 0.235 4.250 ;
    END
END ADDFHX2

MACRO ADDFHX1
    CLASS CORE ;
    FOREIGN ADDFHX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFHXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.945 1.845 14.965 2.075 ;
        RECT  14.715 1.370 14.945 3.520 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.625 1.845 13.645 2.075 ;
        RECT  13.395 1.370 13.625 3.685 ;
        RECT  13.110 3.455 13.395 3.685 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.620 2.940 12.985 3.195 ;
        RECT  12.390 2.350 12.620 3.195 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.905 2.940 7.705 3.375 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.715 1.845 1.105 2.490 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.440 -0.400 15.180 0.400 ;
        RECT  14.100 -0.400 14.440 0.575 ;
        RECT  13.085 -0.400 14.100 0.400 ;
        RECT  12.745 -0.400 13.085 0.575 ;
        RECT  7.655 -0.400 12.745 0.400 ;
        RECT  7.315 -0.400 7.655 0.575 ;
        RECT  1.760 -0.400 7.315 0.400 ;
        RECT  1.420 -0.400 1.760 0.575 ;
        RECT  0.000 -0.400 1.420 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.210 4.640 15.180 5.440 ;
        RECT  13.870 4.465 14.210 5.440 ;
        RECT  11.980 4.640 13.870 5.440 ;
        RECT  11.640 4.465 11.980 5.440 ;
        RECT  7.485 4.640 11.640 5.440 ;
        RECT  7.145 4.065 7.485 5.440 ;
        RECT  2.385 4.640 7.145 5.440 ;
        RECT  2.045 3.690 2.385 5.440 ;
        RECT  1.240 4.640 2.045 5.440 ;
        RECT  0.900 3.755 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.215 2.455 14.305 2.815 ;
        RECT  13.985 2.455 14.215 4.235 ;
        RECT  10.445 4.005 13.985 4.235 ;
        RECT  12.515 0.805 13.790 1.035 ;
        RECT  12.055 1.500 12.915 1.730 ;
        RECT  12.055 3.460 12.745 3.690 ;
        RECT  12.285 0.630 12.515 1.035 ;
        RECT  9.435 0.630 12.285 0.860 ;
        RECT  11.825 1.090 12.055 3.690 ;
        RECT  10.100 1.090 11.825 1.320 ;
        RECT  11.490 2.560 11.825 2.790 ;
        RECT  11.475 1.620 11.595 1.850 ;
        RECT  11.260 1.620 11.475 2.315 ;
        RECT  11.245 1.620 11.260 3.690 ;
        RECT  11.030 2.085 11.245 3.690 ;
        RECT  10.880 3.460 11.030 3.690 ;
        RECT  10.750 1.620 10.875 1.850 ;
        RECT  10.520 1.620 10.750 3.215 ;
        RECT  10.445 2.985 10.520 3.215 ;
        RECT  10.215 2.985 10.445 4.235 ;
        RECT  9.870 1.090 10.100 2.750 ;
        RECT  9.725 2.520 9.870 2.750 ;
        RECT  9.495 2.520 9.725 3.750 ;
        RECT  9.265 0.630 9.435 1.850 ;
        RECT  9.205 0.630 9.265 4.295 ;
        RECT  9.035 1.620 9.205 4.295 ;
        RECT  8.585 4.065 9.035 4.295 ;
        RECT  8.200 0.640 8.905 0.870 ;
        RECT  8.575 1.565 8.805 3.835 ;
        RECT  8.430 1.565 8.575 1.905 ;
        RECT  8.260 3.605 8.575 3.835 ;
        RECT  8.200 2.460 8.345 3.275 ;
        RECT  7.830 3.605 8.260 3.995 ;
        RECT  8.115 0.640 8.200 3.275 ;
        RECT  7.970 0.640 8.115 2.690 ;
        RECT  7.085 0.865 7.970 1.095 ;
        RECT  6.710 3.605 7.830 3.835 ;
        RECT  7.510 1.360 7.740 2.605 ;
        RECT  6.625 1.360 7.510 1.590 ;
        RECT  6.855 0.630 7.085 1.095 ;
        RECT  5.245 0.630 6.855 0.860 ;
        RECT  6.630 3.605 6.710 4.125 ;
        RECT  6.400 2.085 6.630 4.125 ;
        RECT  6.395 1.090 6.625 1.590 ;
        RECT  5.705 1.090 6.395 1.320 ;
        RECT  5.935 1.550 6.165 4.405 ;
        RECT  3.085 4.175 5.935 4.405 ;
        RECT  5.475 1.090 5.705 3.945 ;
        RECT  3.805 3.715 5.475 3.945 ;
        RECT  5.015 0.630 5.245 3.380 ;
        RECT  4.295 0.750 4.525 3.380 ;
        RECT  2.225 0.750 4.295 0.980 ;
        RECT  3.805 1.220 3.860 1.560 ;
        RECT  3.575 1.220 3.805 3.945 ;
        RECT  3.520 1.220 3.575 1.560 ;
        RECT  3.085 1.220 3.140 1.560 ;
        RECT  2.855 1.220 3.085 4.405 ;
        RECT  2.800 1.220 2.855 1.560 ;
        RECT  2.125 2.015 2.605 2.405 ;
        RECT  1.995 0.750 2.225 1.095 ;
        RECT  1.895 1.515 2.125 3.230 ;
        RECT  0.465 0.865 1.995 1.095 ;
        RECT  1.540 1.515 1.895 1.745 ;
        RECT  1.500 3.000 1.895 3.230 ;
        RECT  0.465 3.035 0.520 3.975 ;
        RECT  0.235 0.865 0.465 3.975 ;
        RECT  0.180 3.035 0.235 3.975 ;
    END
END ADDFHX1

MACRO ANTENNA
    CLASS CORE ;
    FOREIGN ANTENNA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.260 0.830 1.780 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.400 1.320 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 4.640 1.320 5.440 ;
        END
    END VDD
END ANTENNA

MACRO RFRDX4
    CLASS CORE ;
    FOREIGN RFRDX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.665 1.460 3.775 1.845 ;
        RECT  3.440 1.460 3.665 2.075 ;
        RECT  3.435 1.460 3.440 2.100 ;
        RECT  3.300 1.845 3.435 2.100 ;
        RECT  3.300 2.635 3.350 3.080 ;
        RECT  3.070 1.845 3.300 3.080 ;
        RECT  1.640 1.845 3.070 2.075 ;
        RECT  3.010 2.635 3.070 3.080 ;
        RECT  1.410 1.845 1.640 2.530 ;
        END
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.410 3.135 2.750 3.475 ;
        RECT  1.535 3.190 2.410 3.420 ;
        RECT  1.355 2.855 1.535 3.420 ;
        RECT  1.180 2.855 1.355 3.760 ;
        RECT  1.180 0.780 1.285 1.615 ;
        RECT  1.175 0.780 1.180 1.845 ;
        RECT  1.175 2.380 1.180 3.780 ;
        RECT  0.945 0.780 1.175 3.780 ;
        RECT  0.800 2.380 0.945 3.780 ;
        END
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 -0.400 3.960 0.400 ;
        RECT  2.010 -0.400 2.045 0.575 ;
        RECT  1.670 -0.400 2.010 1.120 ;
        RECT  0.520 -0.400 1.670 0.400 ;
        RECT  0.520 0.780 0.560 1.120 ;
        RECT  0.220 -0.400 0.520 1.120 ;
        RECT  0.180 -0.400 0.220 0.575 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.160 4.640 3.960 5.440 ;
        RECT  1.820 3.940 2.160 5.440 ;
        RECT  0.560 4.640 1.820 5.440 ;
        RECT  0.220 3.940 0.560 5.440 ;
        RECT  0.000 4.640 0.220 5.440 ;
        END
    END VDD
END RFRDX4

MACRO RFRDX2
    CLASS CORE ;
    FOREIGN RFRDX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RFRDX4 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.030 0.970 3.080 1.310 ;
        RECT  2.800 0.970 3.030 3.655 ;
        RECT  2.740 0.970 2.800 1.310 ;
        RECT  1.105 1.845 2.800 2.075 ;
        RECT  2.690 3.195 2.800 3.655 ;
        RECT  0.875 1.845 1.105 2.600 ;
        END
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 2.785 2.405 3.125 ;
        RECT  1.765 2.840 2.065 3.125 ;
        RECT  0.560 2.840 1.765 3.070 ;
        RECT  0.445 1.460 0.560 1.845 ;
        RECT  0.520 2.840 0.560 3.655 ;
        RECT  0.445 2.635 0.520 3.655 ;
        RECT  0.215 1.460 0.445 3.655 ;
        END
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 -0.400 3.300 0.400 ;
        RECT  1.280 -0.400 1.320 0.575 ;
        RECT  0.940 -0.400 1.280 1.310 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 4.640 3.300 5.440 ;
        RECT  1.020 3.795 1.360 5.440 ;
        RECT  0.000 4.640 1.020 5.440 ;
        END
    END VDD
END RFRDX2

MACRO RFRDX1
    CLASS CORE ;
    FOREIGN RFRDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RFRDX4 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.740 0.970 3.080 1.310 ;
        RECT  2.510 1.080 2.740 1.310 ;
        RECT  2.170 1.080 2.510 3.655 ;
        RECT  2.120 2.075 2.170 2.555 ;
        RECT  1.105 2.325 2.120 2.555 ;
        RECT  0.875 2.200 1.105 2.555 ;
        END
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.855 2.785 1.910 3.125 ;
        RECT  1.570 2.785 1.855 3.195 ;
        RECT  0.560 2.965 1.570 3.195 ;
        RECT  0.330 0.970 0.560 3.655 ;
        RECT  0.220 0.970 0.330 1.310 ;
        RECT  0.220 3.195 0.330 3.655 ;
        END
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 -0.400 3.300 0.400 ;
        RECT  1.280 -0.400 1.320 0.575 ;
        RECT  0.940 -0.400 1.280 1.310 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 4.640 3.300 5.440 ;
        RECT  1.280 4.465 1.320 5.440 ;
        RECT  0.940 3.795 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
END RFRDX1

MACRO XOR3X4
    CLASS CORE ;
    FOREIGN XOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.950 2.940 19.000 4.340 ;
        RECT  18.900 0.955 18.950 4.340 ;
        RECT  18.720 0.835 18.900 4.340 ;
        RECT  18.560 0.835 18.720 1.645 ;
        RECT  18.620 2.740 18.720 4.340 ;
        RECT  18.600 2.740 18.620 3.080 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.350 3.930 17.690 4.270 ;
        RECT  16.945 4.040 17.350 4.270 ;
        RECT  16.715 4.040 16.945 4.315 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.000 2.675 12.110 3.015 ;
        RECT  11.770 1.575 12.000 3.015 ;
        RECT  11.520 1.575 11.770 2.100 ;
        RECT  11.435 1.845 11.520 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.210 1.470 2.550 ;
        RECT  0.875 2.210 1.105 2.635 ;
        RECT  0.660 2.210 0.875 2.550 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 -0.400 19.800 0.400 ;
        RECT  19.280 -0.400 19.620 1.645 ;
        RECT  18.140 -0.400 19.280 0.400 ;
        RECT  17.800 -0.400 18.140 0.630 ;
        RECT  9.375 -0.400 17.800 0.400 ;
        RECT  9.035 -0.400 9.375 0.575 ;
        RECT  7.655 -0.400 9.035 0.400 ;
        RECT  7.315 -0.400 7.655 0.575 ;
        RECT  6.095 -0.400 7.315 0.400 ;
        RECT  5.755 -0.400 6.095 0.575 ;
        RECT  1.280 -0.400 5.755 0.400 ;
        RECT  0.940 -0.400 1.280 1.570 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 4.640 19.800 5.440 ;
        RECT  19.280 3.940 19.620 5.440 ;
        RECT  18.260 4.640 19.280 5.440 ;
        RECT  17.920 3.940 18.260 5.440 ;
        RECT  9.005 4.640 17.920 5.440 ;
        RECT  8.665 4.410 9.005 5.440 ;
        RECT  7.485 4.640 8.665 5.440 ;
        RECT  7.145 4.225 7.485 5.440 ;
        RECT  5.965 4.640 7.145 5.440 ;
        RECT  5.625 4.225 5.965 5.440 ;
        RECT  1.260 4.640 5.625 5.440 ;
        RECT  0.920 3.940 1.260 5.440 ;
        RECT  0.000 4.640 0.920 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.370 2.130 18.490 2.470 ;
        RECT  18.140 2.130 18.370 3.700 ;
        RECT  16.080 3.470 18.140 3.700 ;
        RECT  17.310 1.460 17.540 1.800 ;
        RECT  17.310 2.740 17.500 3.080 ;
        RECT  17.080 1.460 17.310 3.080 ;
        RECT  16.970 2.060 17.080 2.400 ;
        RECT  16.730 0.630 16.840 1.460 ;
        RECT  16.730 2.775 16.800 3.115 ;
        RECT  16.500 0.630 16.730 3.115 ;
        RECT  13.920 0.630 16.500 0.860 ;
        RECT  16.460 2.775 16.500 3.115 ;
        RECT  16.065 1.090 16.120 1.430 ;
        RECT  16.065 2.995 16.080 3.805 ;
        RECT  15.835 1.090 16.065 3.805 ;
        RECT  15.780 1.090 15.835 1.430 ;
        RECT  15.740 2.995 15.835 3.805 ;
        RECT  14.640 1.090 15.780 1.320 ;
        RECT  15.290 1.550 15.400 1.780 ;
        RECT  15.290 2.995 15.360 3.805 ;
        RECT  15.250 1.550 15.290 3.805 ;
        RECT  15.060 1.550 15.250 4.410 ;
        RECT  15.020 2.995 15.060 4.410 ;
        RECT  9.465 4.180 15.020 4.410 ;
        RECT  14.570 1.090 14.640 1.430 ;
        RECT  14.570 2.995 14.640 3.805 ;
        RECT  14.340 1.090 14.570 3.805 ;
        RECT  14.300 1.090 14.340 1.430 ;
        RECT  14.300 2.995 14.340 3.805 ;
        RECT  13.690 0.630 13.920 3.805 ;
        RECT  13.580 0.630 13.690 1.480 ;
        RECT  13.580 2.995 13.690 3.805 ;
        RECT  12.570 0.705 13.580 0.935 ;
        RECT  13.160 3.030 13.200 3.950 ;
        RECT  12.930 1.220 13.160 3.950 ;
        RECT  12.820 1.220 12.930 1.560 ;
        RECT  12.860 3.030 12.930 3.950 ;
        RECT  9.925 3.720 12.860 3.950 ;
        RECT  12.340 0.705 12.570 3.490 ;
        RECT  12.100 1.005 12.340 1.345 ;
        RECT  12.140 3.260 12.340 3.490 ;
        RECT  11.130 1.115 12.100 1.345 ;
        RECT  10.385 3.260 11.675 3.490 ;
        RECT  10.085 0.630 11.530 0.860 ;
        RECT  10.900 1.115 11.130 3.030 ;
        RECT  10.430 1.115 10.900 1.455 ;
        RECT  10.615 2.800 10.900 3.030 ;
        RECT  10.155 2.750 10.385 3.490 ;
        RECT  10.085 2.750 10.155 3.090 ;
        RECT  9.855 0.630 10.085 3.090 ;
        RECT  9.695 3.490 9.925 3.950 ;
        RECT  9.710 0.805 9.855 1.730 ;
        RECT  7.465 0.805 9.710 1.035 ;
        RECT  9.625 3.490 9.695 3.720 ;
        RECT  9.395 2.000 9.625 3.720 ;
        RECT  9.235 3.950 9.465 4.410 ;
        RECT  9.035 2.000 9.395 2.230 ;
        RECT  7.945 3.950 9.235 4.180 ;
        RECT  8.825 2.625 9.165 2.965 ;
        RECT  8.805 1.270 9.035 2.230 ;
        RECT  8.575 2.625 8.825 2.855 ;
        RECT  7.955 1.270 8.805 1.500 ;
        RECT  8.465 1.730 8.575 2.855 ;
        RECT  8.235 1.730 8.465 3.535 ;
        RECT  6.155 3.305 8.235 3.535 ;
        RECT  7.725 1.270 7.955 3.075 ;
        RECT  7.715 3.765 7.945 4.180 ;
        RECT  6.785 2.845 7.725 3.075 ;
        RECT  5.395 3.765 7.715 3.995 ;
        RECT  7.125 0.805 7.465 2.560 ;
        RECT  5.015 0.805 7.125 1.035 ;
        RECT  6.785 1.460 6.895 1.800 ;
        RECT  6.555 1.265 6.785 3.075 ;
        RECT  4.740 1.265 6.555 1.495 ;
        RECT  6.385 2.845 6.555 3.075 ;
        RECT  5.925 1.780 6.155 3.535 ;
        RECT  5.205 1.780 5.925 2.010 ;
        RECT  4.935 3.305 5.925 3.535 ;
        RECT  5.335 2.395 5.445 2.735 ;
        RECT  5.165 3.765 5.395 4.050 ;
        RECT  5.105 2.395 5.335 3.075 ;
        RECT  4.195 3.820 5.165 4.050 ;
        RECT  4.575 2.845 5.105 3.075 ;
        RECT  4.675 0.630 5.015 1.035 ;
        RECT  4.705 3.305 4.935 3.590 ;
        RECT  4.510 1.265 4.740 1.890 ;
        RECT  2.860 3.360 4.705 3.590 ;
        RECT  2.040 0.630 4.675 0.860 ;
        RECT  3.520 1.660 4.510 1.890 ;
        RECT  3.940 1.090 4.280 1.430 ;
        RECT  3.855 3.820 4.195 4.160 ;
        RECT  2.760 1.090 3.940 1.320 ;
        RECT  2.660 3.820 3.855 4.050 ;
        RECT  3.410 1.550 3.520 1.890 ;
        RECT  3.410 2.790 3.435 3.130 ;
        RECT  3.180 1.550 3.410 3.130 ;
        RECT  3.095 2.790 3.180 3.130 ;
        RECT  2.630 2.250 2.860 3.590 ;
        RECT  2.650 1.090 2.760 1.430 ;
        RECT  2.400 3.820 2.660 4.160 ;
        RECT  2.420 1.090 2.650 2.020 ;
        RECT  2.400 1.790 2.420 2.020 ;
        RECT  2.320 1.790 2.400 4.160 ;
        RECT  2.170 1.790 2.320 4.105 ;
        RECT  1.940 0.630 2.040 1.560 ;
        RECT  1.710 0.630 1.940 3.240 ;
        RECT  1.700 0.630 1.710 1.560 ;
        RECT  1.600 2.890 1.710 3.240 ;
        RECT  0.580 2.890 1.600 3.120 ;
        RECT  0.410 2.890 0.580 3.240 ;
        RECT  0.410 0.765 0.520 1.575 ;
        RECT  0.180 0.765 0.410 3.240 ;
    END
END XOR3X4

MACRO XOR3X2
    CLASS CORE ;
    FOREIGN XOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR3X4 ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.700 0.955 11.750 3.025 ;
        RECT  11.665 0.835 11.700 3.080 ;
        RECT  11.520 0.835 11.665 3.195 ;
        RECT  11.360 0.835 11.520 1.645 ;
        RECT  11.435 2.740 11.520 3.195 ;
        RECT  11.360 2.740 11.435 3.080 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.920 3.310 10.450 3.780 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.025 2.405 7.045 2.635 ;
        RECT  6.915 2.405 7.025 3.230 ;
        RECT  6.685 1.790 6.915 3.230 ;
        RECT  6.365 1.790 6.685 2.130 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.210 0.820 2.550 ;
        RECT  0.215 2.210 0.445 2.635 ;
        RECT  0.140 2.210 0.215 2.550 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.940 -0.400 11.880 0.400 ;
        RECT  10.600 -0.400 10.940 0.630 ;
        RECT  3.695 -0.400 10.600 0.400 ;
        RECT  3.355 -0.400 3.695 0.815 ;
        RECT  0.520 -0.400 3.355 0.400 ;
        RECT  0.180 -0.400 0.520 1.570 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.020 4.640 11.880 5.440 ;
        RECT  10.680 3.940 11.020 5.440 ;
        RECT  3.535 4.640 10.680 5.440 ;
        RECT  3.195 4.185 3.535 5.440 ;
        RECT  0.600 4.640 3.195 5.440 ;
        RECT  0.260 3.940 0.600 5.440 ;
        RECT  0.000 4.640 0.260 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.130 2.130 11.290 2.470 ;
        RECT  10.900 1.000 11.130 2.470 ;
        RECT  10.180 1.000 10.900 1.230 ;
        RECT  10.110 1.460 10.340 1.800 ;
        RECT  10.110 2.740 10.300 3.080 ;
        RECT  9.950 0.765 10.180 1.230 ;
        RECT  9.880 1.460 10.110 3.080 ;
        RECT  8.880 0.765 9.950 0.995 ;
        RECT  9.770 2.060 9.880 2.400 ;
        RECT  9.530 1.225 9.640 1.565 ;
        RECT  9.530 2.995 9.600 3.805 ;
        RECT  9.490 1.225 9.530 3.805 ;
        RECT  9.300 1.225 9.490 4.410 ;
        RECT  9.260 2.995 9.300 4.410 ;
        RECT  4.615 4.180 9.260 4.410 ;
        RECT  8.810 0.630 8.880 1.440 ;
        RECT  8.810 2.995 8.880 3.805 ;
        RECT  8.580 0.630 8.810 3.805 ;
        RECT  8.540 0.630 8.580 1.440 ;
        RECT  8.540 2.995 8.580 3.805 ;
        RECT  7.930 0.630 8.160 3.805 ;
        RECT  7.820 0.630 7.930 1.480 ;
        RECT  7.820 2.995 7.930 3.805 ;
        RECT  6.135 0.630 7.820 0.860 ;
        RECT  7.360 1.220 7.590 3.950 ;
        RECT  7.060 1.220 7.360 1.560 ;
        RECT  7.100 3.610 7.360 3.950 ;
        RECT  5.075 3.720 7.100 3.950 ;
        RECT  6.115 2.750 6.455 3.090 ;
        RECT  6.025 0.630 6.135 1.730 ;
        RECT  6.025 2.750 6.115 2.980 ;
        RECT  5.905 0.630 6.025 2.980 ;
        RECT  5.795 0.920 5.905 2.980 ;
        RECT  5.535 3.260 5.735 3.490 ;
        RECT  5.415 1.045 5.535 3.490 ;
        RECT  5.305 0.840 5.415 3.490 ;
        RECT  5.075 0.840 5.305 1.275 ;
        RECT  3.235 1.045 5.075 1.275 ;
        RECT  4.845 1.505 5.075 3.950 ;
        RECT  3.695 1.505 4.845 1.735 ;
        RECT  4.565 1.965 4.615 2.195 ;
        RECT  4.385 3.725 4.615 4.410 ;
        RECT  4.455 1.965 4.565 2.800 ;
        RECT  4.225 1.965 4.455 3.495 ;
        RECT  2.000 3.725 4.385 3.955 ;
        RECT  2.200 3.265 4.225 3.495 ;
        RECT  3.465 1.505 3.695 3.035 ;
        RECT  2.665 2.805 3.465 3.035 ;
        RECT  3.125 1.045 3.235 2.560 ;
        RECT  2.895 0.630 3.125 2.560 ;
        RECT  1.280 0.630 2.895 0.860 ;
        RECT  2.435 1.120 2.665 3.035 ;
        RECT  1.970 2.070 2.200 3.495 ;
        RECT  1.740 1.090 2.000 1.430 ;
        RECT  1.740 3.725 2.000 4.065 ;
        RECT  1.660 1.090 1.740 4.065 ;
        RECT  1.510 1.145 1.660 4.010 ;
        RECT  1.050 0.630 1.280 3.130 ;
        RECT  0.940 0.630 1.050 1.470 ;
        RECT  0.940 2.790 1.050 3.130 ;
    END
END XOR3X2

MACRO XNOR3X4
    CLASS CORE ;
    FOREIGN XNOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.950 2.940 19.000 4.340 ;
        RECT  18.900 0.955 18.950 4.340 ;
        RECT  18.720 0.835 18.900 4.340 ;
        RECT  18.560 0.835 18.720 1.645 ;
        RECT  18.620 2.740 18.720 4.340 ;
        RECT  18.600 2.740 18.620 3.080 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.350 3.930 17.690 4.270 ;
        RECT  16.945 4.040 17.350 4.270 ;
        RECT  16.715 4.040 16.945 4.315 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.960 2.675 12.070 3.015 ;
        RECT  11.730 1.575 11.960 3.015 ;
        RECT  11.520 1.575 11.730 2.100 ;
        RECT  11.435 1.845 11.520 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.210 1.470 2.550 ;
        RECT  0.875 2.210 1.105 2.635 ;
        RECT  0.660 2.210 0.875 2.550 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 -0.400 19.800 0.400 ;
        RECT  19.280 -0.400 19.620 1.645 ;
        RECT  18.140 -0.400 19.280 0.400 ;
        RECT  17.800 -0.400 18.140 0.630 ;
        RECT  9.375 -0.400 17.800 0.400 ;
        RECT  9.035 -0.400 9.375 0.575 ;
        RECT  7.655 -0.400 9.035 0.400 ;
        RECT  7.315 -0.400 7.655 0.575 ;
        RECT  6.095 -0.400 7.315 0.400 ;
        RECT  5.755 -0.400 6.095 0.575 ;
        RECT  1.280 -0.400 5.755 0.400 ;
        RECT  0.940 -0.400 1.280 1.570 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.620 4.640 19.800 5.440 ;
        RECT  19.280 3.940 19.620 5.440 ;
        RECT  18.260 4.640 19.280 5.440 ;
        RECT  17.920 3.940 18.260 5.440 ;
        RECT  9.005 4.640 17.920 5.440 ;
        RECT  8.665 4.410 9.005 5.440 ;
        RECT  7.485 4.640 8.665 5.440 ;
        RECT  7.145 4.225 7.485 5.440 ;
        RECT  5.965 4.640 7.145 5.440 ;
        RECT  5.625 4.225 5.965 5.440 ;
        RECT  1.260 4.640 5.625 5.440 ;
        RECT  0.920 3.940 1.260 5.440 ;
        RECT  0.000 4.640 0.920 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.370 2.130 18.490 2.470 ;
        RECT  18.140 2.130 18.370 3.700 ;
        RECT  16.105 3.470 18.140 3.700 ;
        RECT  17.340 1.460 17.580 1.800 ;
        RECT  17.340 2.740 17.500 3.080 ;
        RECT  17.110 1.460 17.340 3.080 ;
        RECT  16.970 2.095 17.110 2.435 ;
        RECT  16.730 1.460 16.880 1.800 ;
        RECT  16.730 2.775 16.800 3.115 ;
        RECT  16.500 0.630 16.730 3.115 ;
        RECT  13.880 0.630 16.500 0.860 ;
        RECT  16.460 2.775 16.500 3.115 ;
        RECT  16.105 1.090 16.160 1.480 ;
        RECT  16.080 1.090 16.105 3.700 ;
        RECT  15.875 1.090 16.080 3.805 ;
        RECT  15.820 1.090 15.875 1.480 ;
        RECT  15.740 2.995 15.875 3.805 ;
        RECT  14.600 1.090 15.820 1.320 ;
        RECT  15.290 1.550 15.400 1.780 ;
        RECT  15.290 2.995 15.360 3.805 ;
        RECT  15.250 1.550 15.290 3.805 ;
        RECT  15.060 1.550 15.250 4.410 ;
        RECT  15.020 2.995 15.060 4.410 ;
        RECT  9.465 4.180 15.020 4.410 ;
        RECT  14.570 2.995 14.640 3.805 ;
        RECT  14.570 1.090 14.600 1.480 ;
        RECT  14.340 1.090 14.570 3.805 ;
        RECT  14.260 1.090 14.340 1.480 ;
        RECT  14.300 2.995 14.340 3.805 ;
        RECT  13.880 2.995 13.920 3.805 ;
        RECT  13.650 0.630 13.880 3.805 ;
        RECT  13.540 0.630 13.650 1.480 ;
        RECT  13.580 2.995 13.650 3.805 ;
        RECT  12.530 0.705 13.540 0.935 ;
        RECT  13.160 3.030 13.200 3.950 ;
        RECT  12.930 1.220 13.160 3.950 ;
        RECT  12.780 1.220 12.930 1.560 ;
        RECT  12.860 3.030 12.930 3.950 ;
        RECT  9.925 3.720 12.860 3.950 ;
        RECT  12.300 0.705 12.530 3.490 ;
        RECT  12.060 1.005 12.300 1.345 ;
        RECT  12.140 3.260 12.300 3.490 ;
        RECT  11.130 1.115 12.060 1.345 ;
        RECT  10.385 3.260 11.675 3.490 ;
        RECT  10.085 0.630 11.490 0.860 ;
        RECT  10.900 1.115 11.130 3.030 ;
        RECT  10.390 1.115 10.900 1.455 ;
        RECT  10.615 2.800 10.900 3.030 ;
        RECT  10.155 2.745 10.385 3.490 ;
        RECT  10.085 2.745 10.155 3.085 ;
        RECT  9.855 0.630 10.085 3.085 ;
        RECT  9.695 3.490 9.925 3.950 ;
        RECT  9.670 0.805 9.855 1.730 ;
        RECT  9.625 3.490 9.695 3.720 ;
        RECT  7.465 0.805 9.670 1.035 ;
        RECT  9.395 2.000 9.625 3.720 ;
        RECT  9.235 3.950 9.465 4.410 ;
        RECT  9.035 2.000 9.395 2.230 ;
        RECT  7.945 3.950 9.235 4.180 ;
        RECT  8.825 2.625 9.165 2.965 ;
        RECT  8.805 1.270 9.035 2.230 ;
        RECT  8.575 2.625 8.825 2.855 ;
        RECT  7.955 1.270 8.805 1.500 ;
        RECT  8.465 1.730 8.575 2.855 ;
        RECT  8.235 1.730 8.465 3.535 ;
        RECT  6.155 3.305 8.235 3.535 ;
        RECT  7.725 1.270 7.955 3.075 ;
        RECT  7.715 3.765 7.945 4.180 ;
        RECT  6.785 2.845 7.725 3.075 ;
        RECT  5.395 3.765 7.715 3.995 ;
        RECT  7.125 0.805 7.465 2.560 ;
        RECT  5.015 0.805 7.125 1.035 ;
        RECT  6.785 1.460 6.895 1.800 ;
        RECT  6.555 1.265 6.785 3.075 ;
        RECT  4.740 1.265 6.555 1.495 ;
        RECT  6.385 2.845 6.555 3.075 ;
        RECT  5.925 1.725 6.155 3.535 ;
        RECT  5.205 1.725 5.925 2.065 ;
        RECT  4.935 3.305 5.925 3.535 ;
        RECT  5.335 2.395 5.445 2.735 ;
        RECT  5.165 3.765 5.395 4.105 ;
        RECT  5.105 2.395 5.335 3.075 ;
        RECT  4.195 3.875 5.165 4.105 ;
        RECT  4.575 2.845 5.105 3.075 ;
        RECT  4.675 0.630 5.015 1.035 ;
        RECT  4.705 3.305 4.935 3.590 ;
        RECT  4.510 1.265 4.740 1.890 ;
        RECT  2.860 3.360 4.705 3.590 ;
        RECT  2.040 0.630 4.675 0.860 ;
        RECT  3.520 1.660 4.510 1.890 ;
        RECT  3.940 1.090 4.280 1.430 ;
        RECT  3.855 3.820 4.195 4.160 ;
        RECT  2.760 1.090 3.940 1.320 ;
        RECT  2.660 3.820 3.855 4.050 ;
        RECT  3.410 1.550 3.520 1.890 ;
        RECT  3.410 2.790 3.435 3.130 ;
        RECT  3.180 1.550 3.410 3.130 ;
        RECT  3.095 2.790 3.180 3.130 ;
        RECT  2.630 2.250 2.860 3.590 ;
        RECT  2.650 1.090 2.760 1.430 ;
        RECT  2.400 3.820 2.660 4.160 ;
        RECT  2.420 1.090 2.650 2.020 ;
        RECT  2.400 1.790 2.420 2.020 ;
        RECT  2.320 1.790 2.400 4.160 ;
        RECT  2.170 1.790 2.320 4.105 ;
        RECT  1.940 0.630 2.040 1.560 ;
        RECT  1.710 0.630 1.940 3.240 ;
        RECT  1.700 0.630 1.710 1.560 ;
        RECT  1.600 2.890 1.710 3.240 ;
        RECT  0.580 2.890 1.600 3.120 ;
        RECT  0.410 2.890 0.580 3.240 ;
        RECT  0.410 0.765 0.520 1.575 ;
        RECT  0.180 0.765 0.410 3.240 ;
    END
END XNOR3X4

MACRO XNOR3X2
    CLASS CORE ;
    FOREIGN XNOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR3X4 ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.700 0.955 11.750 3.025 ;
        RECT  11.665 0.835 11.700 3.080 ;
        RECT  11.520 0.835 11.665 3.195 ;
        RECT  11.360 0.835 11.520 1.645 ;
        RECT  11.435 2.740 11.520 3.195 ;
        RECT  11.360 2.740 11.435 3.080 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.920 3.310 10.450 3.780 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.025 2.405 7.045 2.635 ;
        RECT  6.915 2.405 7.025 3.230 ;
        RECT  6.685 1.790 6.915 3.230 ;
        RECT  6.365 1.790 6.685 2.130 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.210 0.820 2.550 ;
        RECT  0.215 2.210 0.445 2.635 ;
        RECT  0.140 2.210 0.215 2.550 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.940 -0.400 11.880 0.400 ;
        RECT  10.600 -0.400 10.940 0.630 ;
        RECT  3.695 -0.400 10.600 0.400 ;
        RECT  3.355 -0.400 3.695 0.815 ;
        RECT  0.520 -0.400 3.355 0.400 ;
        RECT  0.180 -0.400 0.520 1.570 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.020 4.640 11.880 5.440 ;
        RECT  10.680 3.940 11.020 5.440 ;
        RECT  3.535 4.640 10.680 5.440 ;
        RECT  3.195 4.185 3.535 5.440 ;
        RECT  0.600 4.640 3.195 5.440 ;
        RECT  0.260 3.940 0.600 5.440 ;
        RECT  0.000 4.640 0.260 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.130 2.130 11.290 2.470 ;
        RECT  10.900 1.000 11.130 2.470 ;
        RECT  10.180 1.000 10.900 1.230 ;
        RECT  10.110 1.460 10.340 1.800 ;
        RECT  10.110 2.740 10.300 3.080 ;
        RECT  9.950 0.630 10.180 1.230 ;
        RECT  9.880 1.460 10.110 3.080 ;
        RECT  8.880 0.630 9.950 0.860 ;
        RECT  9.770 2.210 9.880 2.550 ;
        RECT  9.530 1.140 9.640 1.480 ;
        RECT  9.530 2.995 9.600 3.805 ;
        RECT  9.490 1.140 9.530 3.805 ;
        RECT  9.300 1.140 9.490 4.410 ;
        RECT  9.260 2.995 9.300 4.410 ;
        RECT  4.615 4.180 9.260 4.410 ;
        RECT  8.810 0.630 8.880 1.440 ;
        RECT  8.810 2.995 8.880 3.805 ;
        RECT  8.580 0.630 8.810 3.805 ;
        RECT  8.540 0.630 8.580 1.440 ;
        RECT  8.540 2.995 8.580 3.805 ;
        RECT  7.930 0.630 8.160 3.805 ;
        RECT  7.820 0.630 7.930 1.480 ;
        RECT  7.820 2.995 7.930 3.805 ;
        RECT  6.135 0.630 7.820 0.860 ;
        RECT  7.360 1.220 7.590 3.950 ;
        RECT  7.060 1.220 7.360 1.560 ;
        RECT  7.100 3.610 7.360 3.950 ;
        RECT  5.075 3.720 7.100 3.950 ;
        RECT  6.115 2.750 6.455 3.090 ;
        RECT  6.025 0.630 6.135 1.730 ;
        RECT  6.025 2.750 6.115 2.980 ;
        RECT  5.905 0.630 6.025 2.980 ;
        RECT  5.795 0.920 5.905 2.980 ;
        RECT  5.535 3.260 5.735 3.490 ;
        RECT  5.415 1.045 5.535 3.490 ;
        RECT  5.305 0.840 5.415 3.490 ;
        RECT  5.075 0.840 5.305 1.275 ;
        RECT  3.235 1.045 5.075 1.275 ;
        RECT  4.845 1.505 5.075 3.950 ;
        RECT  3.695 1.505 4.845 1.735 ;
        RECT  4.565 1.965 4.615 2.195 ;
        RECT  4.385 3.725 4.615 4.410 ;
        RECT  4.455 1.965 4.565 2.800 ;
        RECT  4.225 1.965 4.455 3.495 ;
        RECT  2.000 3.725 4.385 3.955 ;
        RECT  2.200 3.265 4.225 3.495 ;
        RECT  3.465 1.505 3.695 3.035 ;
        RECT  2.665 2.805 3.465 3.035 ;
        RECT  3.125 1.045 3.235 2.560 ;
        RECT  2.895 0.630 3.125 2.560 ;
        RECT  1.280 0.630 2.895 0.860 ;
        RECT  2.435 1.120 2.665 3.035 ;
        RECT  1.970 2.070 2.200 3.495 ;
        RECT  1.740 1.090 2.000 1.430 ;
        RECT  1.740 3.725 2.000 4.065 ;
        RECT  1.660 1.090 1.740 4.065 ;
        RECT  1.510 1.145 1.660 4.010 ;
        RECT  1.050 0.630 1.280 3.130 ;
        RECT  0.940 0.630 1.050 1.470 ;
        RECT  0.940 2.790 1.050 3.130 ;
    END
END XNOR3X2

MACRO AFCSHCONX4
    CLASS CORE ;
    FOREIGN AFCSHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 38.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  38.760 0.885 38.800 4.340 ;
        RECT  38.570 0.885 38.760 4.400 ;
        RECT  38.420 0.885 38.570 1.695 ;
        RECT  38.420 2.940 38.570 4.400 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  37.820 1.260 38.140 1.540 ;
        RECT  37.590 1.260 37.820 2.250 ;
        RECT  37.360 2.020 37.590 2.250 ;
        END
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.280 2.175 27.140 2.405 ;
        RECT  24.280 3.615 27.140 3.845 ;
        RECT  23.685 2.175 24.280 3.845 ;
        END
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.125 4.145 21.950 4.375 ;
        RECT  20.170 2.380 20.320 3.780 ;
        RECT  20.125 2.010 20.170 3.780 ;
        RECT  19.940 2.010 20.125 4.375 ;
        RECT  19.350 2.010 19.940 2.240 ;
        RECT  19.895 3.305 19.940 4.375 ;
        RECT  18.400 3.305 19.895 3.535 ;
        END
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  32.690 2.405 32.785 2.635 ;
        RECT  31.935 2.290 32.690 2.635 ;
        RECT  31.410 2.290 31.935 2.630 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.740 2.490 13.545 2.830 ;
        RECT  11.360 2.490 11.740 3.220 ;
        RECT  11.325 2.490 11.360 2.830 ;
        END
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 2.100 5.870 2.820 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 2.180 1.540 2.520 ;
        RECT  0.800 2.180 1.180 3.220 ;
        RECT  0.730 2.180 0.800 2.520 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  38.000 -0.400 38.940 0.400 ;
        RECT  37.660 -0.400 38.000 0.630 ;
        RECT  36.600 -0.400 37.660 0.400 ;
        RECT  36.370 -0.400 36.600 1.750 ;
        RECT  33.500 -0.400 36.370 0.400 ;
        RECT  33.160 -0.400 33.500 0.575 ;
        RECT  31.980 -0.400 33.160 0.400 ;
        RECT  31.640 -0.400 31.980 0.575 ;
        RECT  30.450 -0.400 31.640 0.400 ;
        RECT  30.110 -0.400 30.450 0.575 ;
        RECT  15.300 -0.400 30.110 0.400 ;
        RECT  15.070 -0.400 15.300 0.970 ;
        RECT  13.360 -0.400 15.070 0.400 ;
        RECT  13.020 -0.400 13.360 0.860 ;
        RECT  9.590 -0.400 13.020 0.400 ;
        RECT  8.760 -0.400 9.590 0.960 ;
        RECT  7.575 -0.400 8.760 0.400 ;
        RECT  7.235 -0.400 7.575 0.575 ;
        RECT  6.405 -0.400 7.235 0.400 ;
        RECT  6.065 -0.400 6.405 0.575 ;
        RECT  2.565 -0.400 6.065 0.400 ;
        RECT  2.335 -0.400 2.565 1.020 ;
        RECT  1.360 -0.400 2.335 0.400 ;
        RECT  1.020 -0.400 1.360 1.800 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  38.000 4.640 38.940 5.440 ;
        RECT  37.675 4.465 38.000 5.440 ;
        RECT  37.445 3.665 37.675 5.440 ;
        RECT  36.995 3.665 37.445 3.895 ;
        RECT  33.540 4.640 37.445 5.440 ;
        RECT  33.200 3.450 33.540 5.440 ;
        RECT  31.980 4.640 33.200 5.440 ;
        RECT  31.640 4.465 31.980 5.440 ;
        RECT  30.460 4.640 31.640 5.440 ;
        RECT  30.120 4.465 30.460 5.440 ;
        RECT  14.710 4.640 30.120 5.440 ;
        RECT  14.370 4.465 14.710 5.440 ;
        RECT  13.410 4.640 14.370 5.440 ;
        RECT  13.070 4.465 13.410 5.440 ;
        RECT  11.760 4.640 13.070 5.440 ;
        RECT  11.420 4.465 11.760 5.440 ;
        RECT  10.240 4.640 11.420 5.440 ;
        RECT  9.900 4.465 10.240 5.440 ;
        RECT  8.980 4.640 9.900 5.440 ;
        RECT  8.640 4.465 8.980 5.440 ;
        RECT  6.260 4.640 8.640 5.440 ;
        RECT  5.920 4.465 6.260 5.440 ;
        RECT  2.540 4.640 5.920 5.440 ;
        RECT  2.200 4.090 2.540 5.440 ;
        RECT  1.240 4.640 2.200 5.440 ;
        RECT  0.900 4.090 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  38.190 2.060 38.315 2.710 ;
        RECT  38.085 2.060 38.190 3.435 ;
        RECT  37.960 2.480 38.085 3.435 ;
        RECT  36.765 3.205 37.960 3.435 ;
        RECT  37.110 1.410 37.355 1.750 ;
        RECT  37.110 2.745 37.340 2.975 ;
        RECT  36.880 1.410 37.110 2.975 ;
        RECT  36.305 2.745 36.880 2.975 ;
        RECT  36.535 3.205 36.765 4.405 ;
        RECT  34.925 4.175 36.535 4.405 ;
        RECT  36.075 2.745 36.305 3.915 ;
        RECT  36.140 2.045 36.265 2.275 ;
        RECT  35.910 0.805 36.140 2.275 ;
        RECT  35.385 3.685 36.075 3.915 ;
        RECT  27.730 0.805 35.910 1.035 ;
        RECT  35.680 2.550 35.845 3.450 ;
        RECT  35.615 1.285 35.680 3.450 ;
        RECT  35.450 1.285 35.615 2.780 ;
        RECT  35.185 3.010 35.385 3.915 ;
        RECT  35.155 2.170 35.185 3.915 ;
        RECT  34.955 2.170 35.155 3.240 ;
        RECT  34.720 1.380 35.015 1.720 ;
        RECT  34.720 3.470 34.925 4.405 ;
        RECT  34.695 1.380 34.720 4.405 ;
        RECT  34.490 1.380 34.695 3.770 ;
        RECT  34.205 1.360 34.240 3.340 ;
        RECT  34.010 1.360 34.205 3.965 ;
        RECT  33.975 3.110 34.010 3.965 ;
        RECT  33.550 1.265 33.780 2.670 ;
        RECT  29.120 1.265 33.550 1.495 ;
        RECT  33.090 1.725 33.320 3.130 ;
        RECT  32.400 1.725 33.090 1.955 ;
        RECT  32.765 2.900 33.090 3.130 ;
        RECT  32.535 2.900 32.765 4.280 ;
        RECT  27.660 4.000 32.535 4.230 ;
        RECT  31.165 1.725 31.220 1.955 ;
        RECT  30.860 1.725 31.165 3.770 ;
        RECT  30.855 2.510 30.860 3.770 ;
        RECT  30.075 2.510 30.855 2.740 ;
        RECT  28.420 3.540 30.855 3.770 ;
        RECT  29.845 2.380 30.075 2.740 ;
        RECT  29.610 3.080 29.900 3.310 ;
        RECT  29.610 1.725 29.730 1.955 ;
        RECT  29.380 1.725 29.610 3.310 ;
        RECT  29.350 1.725 29.380 1.955 ;
        RECT  29.120 2.770 29.125 3.310 ;
        RECT  28.895 1.265 29.120 3.310 ;
        RECT  28.890 1.265 28.895 3.000 ;
        RECT  28.630 1.575 28.890 1.805 ;
        RECT  28.195 3.280 28.420 3.770 ;
        RECT  28.080 1.370 28.195 3.770 ;
        RECT  27.965 1.370 28.080 3.510 ;
        RECT  27.500 0.805 27.730 1.945 ;
        RECT  27.430 2.895 27.660 4.230 ;
        RECT  23.405 1.715 27.500 1.945 ;
        RECT  24.565 2.895 27.430 3.125 ;
        RECT  22.810 0.735 27.260 0.965 ;
        RECT  22.055 1.255 27.140 1.485 ;
        RECT  23.175 1.715 23.405 3.915 ;
        RECT  20.780 3.685 23.175 3.915 ;
        RECT  22.385 2.165 22.615 3.455 ;
        RECT  21.490 2.165 22.385 2.395 ;
        RECT  21.010 3.225 22.385 3.455 ;
        RECT  21.825 0.630 22.055 1.485 ;
        RECT  15.760 0.630 21.825 0.860 ;
        RECT  21.260 1.090 21.490 2.395 ;
        RECT  16.220 1.090 21.260 1.320 ;
        RECT  20.550 1.550 20.780 3.915 ;
        RECT  17.250 1.550 20.550 1.780 ;
        RECT  18.170 3.765 19.460 3.995 ;
        RECT  18.860 2.010 18.970 2.240 ;
        RECT  18.630 2.010 18.860 2.745 ;
        RECT  18.170 2.515 18.630 2.745 ;
        RECT  17.710 2.010 18.270 2.240 ;
        RECT  17.940 2.515 18.170 4.235 ;
        RECT  3.145 4.005 17.940 4.235 ;
        RECT  17.480 2.010 17.710 3.270 ;
        RECT  17.470 3.040 17.480 3.270 ;
        RECT  17.240 3.040 17.470 3.775 ;
        RECT  17.020 1.550 17.250 2.810 ;
        RECT  14.935 3.545 17.240 3.775 ;
        RECT  17.010 2.580 17.020 2.810 ;
        RECT  16.780 2.580 17.010 3.315 ;
        RECT  16.680 1.550 16.790 1.780 ;
        RECT  16.135 3.085 16.780 3.315 ;
        RECT  16.550 1.550 16.680 2.350 ;
        RECT  16.450 1.550 16.550 2.810 ;
        RECT  16.320 2.120 16.450 2.810 ;
        RECT  15.755 2.580 16.320 2.810 ;
        RECT  15.990 1.090 16.220 1.890 ;
        RECT  15.200 2.120 16.090 2.350 ;
        RECT  14.740 1.660 15.990 1.890 ;
        RECT  15.530 0.630 15.760 1.430 ;
        RECT  15.525 2.580 15.755 3.315 ;
        RECT  14.280 1.200 15.530 1.430 ;
        RECT  15.410 3.085 15.525 3.315 ;
        RECT  14.970 2.120 15.200 2.870 ;
        RECT  14.935 2.640 14.970 2.870 ;
        RECT  14.705 2.640 14.935 3.775 ;
        RECT  13.820 0.740 14.740 0.970 ;
        RECT  14.510 1.660 14.740 2.260 ;
        RECT  11.000 3.545 14.705 3.775 ;
        RECT  14.290 2.030 14.510 2.260 ;
        RECT  14.060 2.030 14.290 3.310 ;
        RECT  14.050 1.200 14.280 1.780 ;
        RECT  11.870 2.030 14.060 2.260 ;
        RECT  12.250 3.080 14.060 3.310 ;
        RECT  12.330 1.550 14.050 1.780 ;
        RECT  13.590 0.740 13.820 1.320 ;
        RECT  12.790 1.090 13.590 1.320 ;
        RECT  12.560 0.630 12.790 1.320 ;
        RECT  10.145 0.630 12.560 0.860 ;
        RECT  12.100 1.200 12.330 1.780 ;
        RECT  10.610 1.200 12.100 1.430 ;
        RECT  11.460 1.660 11.870 2.260 ;
        RECT  10.775 3.435 11.000 3.775 ;
        RECT  10.660 2.110 10.775 3.775 ;
        RECT  10.545 2.110 10.660 3.720 ;
        RECT  10.380 1.200 10.610 1.880 ;
        RECT  10.200 2.110 10.545 2.340 ;
        RECT  9.480 3.490 10.545 3.720 ;
        RECT  7.145 1.650 10.380 1.880 ;
        RECT  9.915 0.630 10.145 1.420 ;
        RECT  8.030 1.190 9.915 1.420 ;
        RECT  9.140 3.435 9.480 3.775 ;
        RECT  7.955 3.545 8.140 3.775 ;
        RECT  7.800 0.885 8.030 1.420 ;
        RECT  7.725 3.085 7.955 3.775 ;
        RECT  6.380 0.885 7.800 1.115 ;
        RECT  6.380 3.085 7.725 3.315 ;
        RECT  3.980 3.545 7.495 3.775 ;
        RECT  7.145 2.625 7.485 2.855 ;
        RECT  6.915 1.345 7.145 2.855 ;
        RECT  6.810 1.345 6.915 1.880 ;
        RECT  6.625 1.345 6.810 1.575 ;
        RECT  6.150 0.885 6.380 3.315 ;
        RECT  5.125 1.515 5.645 1.745 ;
        RECT  5.160 3.085 5.500 3.315 ;
        RECT  5.125 2.370 5.160 3.315 ;
        RECT  4.930 1.515 5.125 3.315 ;
        RECT  4.765 0.760 5.105 1.100 ;
        RECT  4.895 1.515 4.930 2.600 ;
        RECT  4.665 0.815 4.765 1.100 ;
        RECT  4.665 2.970 4.700 3.310 ;
        RECT  4.435 0.815 4.665 3.310 ;
        RECT  3.025 0.815 4.435 1.045 ;
        RECT  4.360 2.970 4.435 3.310 ;
        RECT  4.030 1.450 4.205 2.605 ;
        RECT  3.980 1.450 4.030 3.145 ;
        RECT  3.975 1.450 3.980 3.775 ;
        RECT  3.800 2.375 3.975 3.775 ;
        RECT  3.640 2.915 3.800 3.775 ;
        RECT  3.260 1.460 3.485 2.455 ;
        RECT  3.255 1.460 3.260 3.305 ;
        RECT  3.030 2.225 3.255 3.305 ;
        RECT  2.915 3.595 3.145 4.235 ;
        RECT  2.920 2.965 3.030 3.305 ;
        RECT  2.795 0.815 3.025 1.480 ;
        RECT  0.520 3.595 2.915 3.825 ;
        RECT  2.080 1.250 2.795 1.480 ;
        RECT  2.080 2.110 2.780 2.450 ;
        RECT  1.960 1.250 2.080 3.070 ;
        RECT  1.850 1.250 1.960 3.180 ;
        RECT  1.740 1.460 1.850 1.800 ;
        RECT  1.620 2.840 1.850 3.180 ;
        RECT  0.410 0.680 0.640 1.800 ;
        RECT  0.410 2.875 0.520 4.155 ;
        RECT  0.300 0.680 0.410 4.155 ;
        RECT  0.180 1.125 0.300 4.155 ;
    END
END AFCSHCONX4

MACRO AFCSHCONX2
    CLASS CORE ;
    FOREIGN AFCSHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFCSHCONX4 ;
    SIZE 33.660 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  33.480 0.885 33.520 4.340 ;
        RECT  33.290 0.885 33.480 4.400 ;
        RECT  33.140 0.885 33.290 1.695 ;
        RECT  33.140 2.940 33.290 4.400 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  32.540 1.260 32.860 1.540 ;
        RECT  32.310 1.260 32.540 2.250 ;
        RECT  32.080 2.020 32.310 2.250 ;
        END
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.690 2.175 22.760 2.405 ;
        RECT  19.690 3.615 20.690 3.845 ;
        RECT  19.460 2.175 19.690 3.845 ;
        RECT  19.280 2.175 19.460 3.220 ;
        END
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.000 3.505 19.230 4.410 ;
        RECT  17.275 4.180 19.000 4.410 ;
        RECT  17.045 3.305 17.275 4.410 ;
        RECT  17.020 3.305 17.045 3.535 ;
        RECT  16.870 2.380 17.020 3.535 ;
        RECT  16.640 2.010 16.870 3.535 ;
        RECT  16.500 2.010 16.640 2.240 ;
        RECT  15.550 3.305 16.640 3.535 ;
        END
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.950 2.230 27.505 2.635 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.420 2.405 10.820 2.745 ;
        RECT  10.040 2.405 10.420 3.220 ;
        RECT  10.010 2.405 10.040 2.745 ;
        END
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.280 2.270 5.800 2.820 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 2.175 1.180 3.220 ;
        RECT  0.800 2.380 0.840 3.220 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  32.720 -0.400 33.660 0.400 ;
        RECT  32.380 -0.400 32.720 0.630 ;
        RECT  31.320 -0.400 32.380 0.400 ;
        RECT  31.090 -0.400 31.320 1.750 ;
        RECT  28.220 -0.400 31.090 0.400 ;
        RECT  27.880 -0.400 28.220 0.575 ;
        RECT  25.990 -0.400 27.880 0.400 ;
        RECT  25.650 -0.400 25.990 0.575 ;
        RECT  12.450 -0.400 25.650 0.400 ;
        RECT  12.220 -0.400 12.450 0.970 ;
        RECT  8.945 -0.400 12.220 0.400 ;
        RECT  8.605 -0.400 8.945 0.960 ;
        RECT  7.425 -0.400 8.605 0.400 ;
        RECT  7.085 -0.400 7.425 0.575 ;
        RECT  6.060 -0.400 7.085 0.400 ;
        RECT  5.720 -0.400 6.060 0.575 ;
        RECT  2.500 -0.400 5.720 0.400 ;
        RECT  2.160 -0.400 2.500 0.575 ;
        RECT  1.200 -0.400 2.160 0.400 ;
        RECT  0.860 -0.400 1.200 0.575 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  32.720 4.640 33.660 5.440 ;
        RECT  32.380 4.465 32.720 5.440 ;
        RECT  32.105 4.640 32.380 5.440 ;
        RECT  31.875 3.665 32.105 5.440 ;
        RECT  31.715 3.665 31.875 3.895 ;
        RECT  28.260 4.640 31.875 5.440 ;
        RECT  27.920 3.450 28.260 5.440 ;
        RECT  26.080 4.640 27.920 5.440 ;
        RECT  25.740 4.465 26.080 5.440 ;
        RECT  11.860 4.640 25.740 5.440 ;
        RECT  11.520 4.465 11.860 5.440 ;
        RECT  10.200 4.640 11.520 5.440 ;
        RECT  9.860 4.465 10.200 5.440 ;
        RECT  8.680 4.640 9.860 5.440 ;
        RECT  8.340 4.465 8.680 5.440 ;
        RECT  6.140 4.640 8.340 5.440 ;
        RECT  5.800 4.465 6.140 5.440 ;
        RECT  2.420 4.640 5.800 5.440 ;
        RECT  2.080 4.465 2.420 5.440 ;
        RECT  1.160 4.640 2.080 5.440 ;
        RECT  0.820 4.090 1.160 5.440 ;
        RECT  0.000 4.640 0.820 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  32.910 2.060 33.035 2.710 ;
        RECT  32.805 2.060 32.910 3.435 ;
        RECT  32.680 2.480 32.805 3.435 ;
        RECT  31.485 3.205 32.680 3.435 ;
        RECT  31.830 1.410 32.075 1.750 ;
        RECT  31.830 2.745 32.060 2.975 ;
        RECT  31.600 1.410 31.830 2.975 ;
        RECT  31.025 2.745 31.600 2.975 ;
        RECT  31.255 3.205 31.485 4.405 ;
        RECT  29.645 4.175 31.255 4.405 ;
        RECT  30.795 2.745 31.025 3.915 ;
        RECT  30.860 2.045 30.985 2.275 ;
        RECT  30.630 0.805 30.860 2.275 ;
        RECT  30.105 3.685 30.795 3.915 ;
        RECT  23.270 0.805 30.630 1.035 ;
        RECT  30.400 2.505 30.565 3.450 ;
        RECT  30.335 1.285 30.400 3.450 ;
        RECT  30.170 1.285 30.335 2.735 ;
        RECT  29.905 2.965 30.105 3.915 ;
        RECT  29.875 2.170 29.905 3.915 ;
        RECT  29.675 2.170 29.875 3.195 ;
        RECT  29.440 1.380 29.735 1.720 ;
        RECT  29.440 3.425 29.645 4.405 ;
        RECT  29.415 1.380 29.440 4.405 ;
        RECT  29.210 1.380 29.415 3.655 ;
        RECT  28.925 1.360 28.960 3.130 ;
        RECT  28.730 1.360 28.925 4.260 ;
        RECT  28.695 2.900 28.730 4.260 ;
        RECT  28.270 1.265 28.500 2.670 ;
        RECT  24.660 1.265 28.270 1.495 ;
        RECT  27.810 1.725 28.040 3.130 ;
        RECT  27.120 1.725 27.810 1.955 ;
        RECT  27.485 2.900 27.810 3.130 ;
        RECT  27.255 2.900 27.485 4.280 ;
        RECT  22.825 4.000 27.255 4.230 ;
        RECT  26.705 2.960 26.785 3.770 ;
        RECT  26.705 1.725 26.760 1.955 ;
        RECT  26.475 1.725 26.705 3.770 ;
        RECT  26.400 1.725 26.475 2.770 ;
        RECT  24.040 3.540 26.475 3.770 ;
        RECT  25.695 2.510 26.400 2.740 ;
        RECT  25.465 2.380 25.695 2.740 ;
        RECT  25.210 3.080 25.520 3.310 ;
        RECT  25.210 1.725 25.270 1.955 ;
        RECT  24.980 1.725 25.210 3.310 ;
        RECT  24.890 1.725 24.980 1.955 ;
        RECT  24.660 2.770 24.745 3.310 ;
        RECT  24.515 1.265 24.660 3.310 ;
        RECT  24.430 1.265 24.515 3.000 ;
        RECT  24.170 1.575 24.430 1.805 ;
        RECT  23.735 3.280 24.040 3.770 ;
        RECT  23.700 1.370 23.735 3.770 ;
        RECT  23.505 1.370 23.700 3.510 ;
        RECT  23.040 0.805 23.270 1.945 ;
        RECT  18.770 1.715 23.040 1.945 ;
        RECT  22.595 2.895 22.825 4.230 ;
        RECT  18.630 0.735 22.810 0.965 ;
        RECT  18.400 1.255 22.760 1.485 ;
        RECT  20.125 2.895 22.595 3.125 ;
        RECT  18.540 1.715 18.770 3.950 ;
        RECT  17.735 3.720 18.540 3.950 ;
        RECT  18.170 0.630 18.400 1.485 ;
        RECT  18.080 2.165 18.310 3.490 ;
        RECT  12.910 0.630 18.170 0.860 ;
        RECT  17.940 2.165 18.080 2.395 ;
        RECT  17.965 3.260 18.080 3.490 ;
        RECT  17.710 1.090 17.940 2.395 ;
        RECT  17.505 2.675 17.735 3.950 ;
        RECT  13.370 1.090 17.710 1.320 ;
        RECT  17.480 2.675 17.505 2.905 ;
        RECT  17.250 1.550 17.480 2.905 ;
        RECT  14.400 1.550 17.250 1.780 ;
        RECT  15.320 3.765 16.610 3.995 ;
        RECT  16.010 2.010 16.120 2.240 ;
        RECT  15.780 2.010 16.010 2.745 ;
        RECT  15.320 2.515 15.780 2.745 ;
        RECT  14.860 2.010 15.420 2.240 ;
        RECT  15.090 2.515 15.320 4.235 ;
        RECT  3.170 4.005 15.090 4.235 ;
        RECT  14.630 2.010 14.860 3.270 ;
        RECT  14.620 3.040 14.630 3.270 ;
        RECT  14.390 3.040 14.620 3.775 ;
        RECT  14.170 1.550 14.400 2.810 ;
        RECT  12.085 3.545 14.390 3.775 ;
        RECT  14.160 2.580 14.170 2.810 ;
        RECT  13.930 2.580 14.160 3.315 ;
        RECT  13.830 1.550 13.940 1.780 ;
        RECT  13.285 3.085 13.930 3.315 ;
        RECT  13.700 1.550 13.830 2.350 ;
        RECT  13.600 1.550 13.700 2.810 ;
        RECT  13.470 2.120 13.600 2.810 ;
        RECT  12.905 2.580 13.470 2.810 ;
        RECT  13.140 1.090 13.370 1.890 ;
        RECT  12.085 2.120 13.240 2.350 ;
        RECT  11.280 1.660 13.140 1.890 ;
        RECT  12.680 0.630 12.910 1.430 ;
        RECT  12.675 2.580 12.905 3.315 ;
        RECT  9.920 1.200 12.680 1.430 ;
        RECT  12.560 3.085 12.675 3.315 ;
        RECT  11.855 2.120 12.085 3.775 ;
        RECT  9.455 0.735 11.890 0.965 ;
        RECT  9.775 3.545 11.855 3.775 ;
        RECT  11.050 1.660 11.280 3.310 ;
        RECT  11.020 1.660 11.050 1.890 ;
        RECT  10.700 3.080 11.050 3.310 ;
        RECT  9.690 1.200 9.920 1.880 ;
        RECT  9.545 2.110 9.775 3.775 ;
        RECT  7.000 1.650 9.690 1.880 ;
        RECT  9.420 2.110 9.545 2.340 ;
        RECT  9.100 3.435 9.545 3.775 ;
        RECT  9.225 0.735 9.455 1.420 ;
        RECT  7.795 1.190 9.225 1.420 ;
        RECT  7.810 3.370 7.920 3.710 ;
        RECT  7.580 3.085 7.810 3.710 ;
        RECT  7.565 0.875 7.795 1.420 ;
        RECT  6.260 3.085 7.580 3.315 ;
        RECT  6.085 0.875 7.565 1.105 ;
        RECT  3.860 3.545 7.270 3.775 ;
        RECT  7.000 2.625 7.140 2.855 ;
        RECT  6.770 1.345 7.000 2.855 ;
        RECT  6.480 1.345 6.770 1.575 ;
        RECT  6.085 1.805 6.260 3.315 ;
        RECT  6.030 0.875 6.085 3.315 ;
        RECT  5.855 0.875 6.030 2.035 ;
        RECT  5.040 3.085 5.380 3.315 ;
        RECT  4.945 1.515 5.290 1.745 ;
        RECT  4.945 2.290 5.040 3.315 ;
        RECT  4.810 1.515 4.945 3.315 ;
        RECT  4.715 1.515 4.810 2.520 ;
        RECT  4.475 0.760 4.760 1.165 ;
        RECT  4.475 2.970 4.580 3.310 ;
        RECT  4.420 0.760 4.475 3.310 ;
        RECT  4.245 0.935 4.420 3.310 ;
        RECT  1.880 0.935 4.245 1.165 ;
        RECT  4.240 2.970 4.245 3.310 ;
        RECT  3.805 1.450 3.980 1.790 ;
        RECT  3.805 2.965 3.860 3.775 ;
        RECT  3.575 1.450 3.805 3.775 ;
        RECT  3.520 2.965 3.575 3.775 ;
        RECT  3.100 1.460 3.260 1.800 ;
        RECT  2.940 3.570 3.170 4.235 ;
        RECT  2.870 1.460 3.100 3.110 ;
        RECT  0.520 3.570 2.940 3.800 ;
        RECT  2.760 2.770 2.870 3.110 ;
        RECT  1.880 2.110 2.585 2.450 ;
        RECT  1.650 0.935 1.880 3.080 ;
        RECT  1.540 1.460 1.650 1.800 ;
        RECT  1.460 2.740 1.650 3.080 ;
        RECT  0.290 1.460 0.520 3.800 ;
        RECT  0.180 1.460 0.290 1.800 ;
        RECT  0.180 2.810 0.290 3.150 ;
    END
END AFCSHCONX2

MACRO AFCSHCINX4
    CLASS CORE ;
    FOREIGN AFCSHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 38.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  37.910 0.990 38.140 4.340 ;
        RECT  37.760 0.990 37.910 1.800 ;
        RECT  37.760 2.940 37.910 4.340 ;
        RECT  37.650 2.940 37.760 4.220 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  37.175 1.285 37.405 1.540 ;
        RECT  36.895 1.310 37.175 1.540 ;
        RECT  36.665 1.310 36.895 2.460 ;
        END
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  25.560 2.155 26.370 2.495 ;
        RECT  25.405 3.595 26.215 3.935 ;
        RECT  25.155 2.155 25.560 2.385 ;
        RECT  24.635 3.595 25.405 3.825 ;
        RECT  24.925 1.730 25.155 2.385 ;
        RECT  24.865 1.730 24.925 2.075 ;
        RECT  23.025 1.730 24.865 1.960 ;
        RECT  24.405 3.260 24.635 3.825 ;
        RECT  23.025 3.260 24.405 3.490 ;
        RECT  22.795 1.730 23.025 3.490 ;
        RECT  22.580 1.820 22.795 3.220 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.640 1.870 21.870 3.490 ;
        RECT  20.980 1.870 21.640 2.100 ;
        RECT  17.480 3.260 21.640 3.490 ;
        RECT  20.650 1.260 20.980 2.100 ;
        RECT  20.600 1.260 20.650 2.570 ;
        RECT  20.420 1.870 20.600 2.570 ;
        RECT  18.595 2.340 20.420 2.570 ;
        RECT  18.365 1.820 18.595 2.570 ;
        RECT  18.265 1.820 18.365 2.100 ;
        RECT  17.400 1.820 18.265 2.050 ;
        END
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  31.495 2.270 32.170 2.755 ;
        RECT  31.320 2.320 31.495 2.660 ;
        END
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 2.055 10.050 2.660 ;
        END
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 2.245 8.685 2.700 ;
        RECT  7.860 2.470 8.060 2.700 ;
        RECT  7.630 2.470 7.860 3.315 ;
        RECT  6.595 3.085 7.630 3.315 ;
        RECT  6.365 1.390 6.595 3.315 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.490 2.105 1.600 2.445 ;
        RECT  1.260 2.105 1.490 2.850 ;
        RECT  1.180 2.620 1.260 2.850 ;
        RECT  0.950 2.620 1.180 3.195 ;
        RECT  0.875 2.965 0.950 3.195 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  37.335 -0.400 38.280 0.400 ;
        RECT  36.995 -0.400 37.335 0.575 ;
        RECT  35.960 -0.400 36.995 0.400 ;
        RECT  35.620 -0.400 35.960 1.100 ;
        RECT  32.585 -0.400 35.620 0.400 ;
        RECT  32.245 -0.400 32.585 0.575 ;
        RECT  31.065 -0.400 32.245 0.400 ;
        RECT  30.725 -0.400 31.065 0.575 ;
        RECT  29.965 -0.400 30.725 0.400 ;
        RECT  29.625 -0.400 29.965 0.575 ;
        RECT  13.480 -0.400 29.625 0.400 ;
        RECT  12.200 -0.400 13.480 0.575 ;
        RECT  7.610 -0.400 12.200 0.400 ;
        RECT  6.800 -0.400 7.610 0.575 ;
        RECT  2.400 -0.400 6.800 0.400 ;
        RECT  2.060 -0.400 2.400 0.575 ;
        RECT  1.280 -0.400 2.060 0.400 ;
        RECT  0.940 -0.400 1.280 0.630 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  37.230 4.640 38.280 5.440 ;
        RECT  36.890 3.830 37.230 5.440 ;
        RECT  36.420 4.640 36.890 5.440 ;
        RECT  36.080 3.760 36.420 5.440 ;
        RECT  32.610 4.640 36.080 5.440 ;
        RECT  32.270 3.150 32.610 5.440 ;
        RECT  31.130 4.640 32.270 5.440 ;
        RECT  30.790 4.465 31.130 5.440 ;
        RECT  30.015 4.640 30.790 5.440 ;
        RECT  29.675 4.465 30.015 5.440 ;
        RECT  10.335 4.640 29.675 5.440 ;
        RECT  9.055 4.465 10.335 5.440 ;
        RECT  8.090 4.640 9.055 5.440 ;
        RECT  7.750 4.465 8.090 5.440 ;
        RECT  2.390 4.640 7.750 5.440 ;
        RECT  2.050 4.465 2.390 5.440 ;
        RECT  1.240 4.640 2.050 5.440 ;
        RECT  0.900 4.080 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  37.410 2.170 37.680 2.535 ;
        RECT  37.340 2.170 37.410 3.530 ;
        RECT  37.180 2.305 37.340 3.530 ;
        RECT  35.850 3.300 37.180 3.530 ;
        RECT  36.325 2.840 36.470 3.070 ;
        RECT  36.325 1.460 36.435 1.800 ;
        RECT  36.095 1.460 36.325 3.070 ;
        RECT  35.390 2.840 36.095 3.070 ;
        RECT  35.620 3.300 35.850 4.405 ;
        RECT  34.010 4.175 35.620 4.405 ;
        RECT  35.390 2.100 35.500 2.440 ;
        RECT  35.160 0.805 35.390 2.440 ;
        RECT  35.160 2.840 35.390 3.915 ;
        RECT  29.055 0.805 35.160 1.035 ;
        RECT  34.470 3.685 35.160 3.915 ;
        RECT  34.700 1.380 34.930 3.450 ;
        RECT  34.445 1.380 34.700 1.720 ;
        RECT  34.240 2.170 34.470 3.915 ;
        RECT  34.010 1.380 34.065 1.720 ;
        RECT  33.780 1.380 34.010 4.405 ;
        RECT  33.725 1.380 33.780 1.720 ;
        RECT  33.275 1.460 33.345 1.800 ;
        RECT  33.275 3.110 33.345 4.390 ;
        RECT  33.045 1.460 33.275 4.390 ;
        RECT  33.005 1.460 33.045 1.800 ;
        RECT  33.005 3.110 33.045 4.390 ;
        RECT  32.690 2.440 32.800 2.780 ;
        RECT  32.460 1.265 32.690 2.780 ;
        RECT  28.370 1.265 32.460 1.495 ;
        RECT  31.550 3.110 31.890 4.390 ;
        RECT  31.090 1.730 31.825 1.960 ;
        RECT  31.090 3.720 31.550 3.950 ;
        RECT  30.860 1.730 31.090 3.950 ;
        RECT  27.860 3.720 30.860 3.950 ;
        RECT  30.285 1.730 30.515 3.310 ;
        RECT  30.125 1.730 30.285 2.565 ;
        RECT  29.215 2.335 30.125 2.565 ;
        RECT  28.985 2.965 29.190 3.305 ;
        RECT  28.985 1.725 29.185 1.955 ;
        RECT  28.825 0.635 29.055 1.035 ;
        RECT  28.755 1.725 28.985 3.305 ;
        RECT  11.200 4.180 28.895 4.410 ;
        RECT  20.185 0.635 28.825 0.865 ;
        RECT  28.370 3.150 28.525 3.490 ;
        RECT  28.140 1.265 28.370 3.490 ;
        RECT  27.630 1.335 27.860 3.950 ;
        RECT  27.365 1.335 27.630 1.675 ;
        RECT  27.465 2.985 27.630 3.950 ;
        RECT  26.330 2.985 27.465 3.215 ;
        RECT  25.790 1.375 26.370 1.715 ;
        RECT  25.750 2.875 26.330 3.215 ;
        RECT  25.560 1.180 25.790 1.715 ;
        RECT  25.520 2.790 25.750 3.215 ;
        RECT  22.350 1.180 25.560 1.410 ;
        RECT  23.745 2.790 25.520 3.020 ;
        RECT  23.405 2.210 23.745 3.020 ;
        RECT  22.120 1.180 22.350 3.950 ;
        RECT  21.965 1.180 22.120 1.410 ;
        RECT  11.660 3.720 22.120 3.950 ;
        RECT  20.920 2.685 21.150 3.030 ;
        RECT  18.135 2.800 20.920 3.030 ;
        RECT  19.955 0.635 20.185 2.110 ;
        RECT  19.055 1.880 19.955 2.110 ;
        RECT  19.515 1.420 19.725 1.650 ;
        RECT  19.285 0.840 19.515 1.650 ;
        RECT  17.865 0.840 19.285 1.070 ;
        RECT  18.825 1.350 19.055 2.110 ;
        RECT  17.330 1.350 18.825 1.580 ;
        RECT  17.905 2.485 18.135 3.030 ;
        RECT  17.325 2.485 17.905 2.825 ;
        RECT  17.635 0.630 17.865 1.070 ;
        RECT  14.675 0.630 17.635 0.860 ;
        RECT  17.100 1.090 17.330 1.580 ;
        RECT  16.710 2.540 17.325 2.770 ;
        RECT  15.995 1.090 17.100 1.320 ;
        RECT  16.710 1.550 16.865 1.780 ;
        RECT  16.480 1.550 16.710 3.490 ;
        RECT  12.120 3.260 16.480 3.490 ;
        RECT  15.885 1.090 15.995 1.525 ;
        RECT  15.655 1.090 15.885 3.030 ;
        RECT  15.240 2.800 15.655 3.030 ;
        RECT  14.995 1.190 15.135 2.060 ;
        RECT  14.905 1.190 14.995 3.030 ;
        RECT  14.765 1.830 14.905 3.030 ;
        RECT  14.520 2.800 14.765 3.030 ;
        RECT  14.445 0.630 14.675 1.495 ;
        RECT  11.500 1.265 14.445 1.495 ;
        RECT  14.025 2.385 14.255 3.030 ;
        RECT  14.020 0.630 14.215 0.860 ;
        RECT  12.580 2.800 14.025 3.030 ;
        RECT  13.790 0.630 14.020 1.035 ;
        RECT  11.960 0.805 13.790 1.035 ;
        RECT  12.350 1.725 12.580 3.030 ;
        RECT  11.960 1.725 12.350 1.955 ;
        RECT  11.890 3.085 12.120 3.490 ;
        RECT  11.730 0.630 11.960 1.035 ;
        RECT  10.985 3.085 11.890 3.315 ;
        RECT  8.070 0.630 11.730 0.860 ;
        RECT  11.430 3.545 11.660 3.950 ;
        RECT  11.270 1.090 11.500 1.495 ;
        RECT  6.595 3.545 11.430 3.775 ;
        RECT  8.530 1.090 11.270 1.320 ;
        RECT  10.970 4.005 11.200 4.410 ;
        RECT  10.985 1.550 11.040 1.890 ;
        RECT  10.755 1.550 10.985 3.315 ;
        RECT  7.270 4.005 10.970 4.235 ;
        RECT  10.700 1.550 10.755 1.890 ;
        RECT  9.815 3.085 10.755 3.315 ;
        RECT  8.920 1.550 9.150 3.205 ;
        RECT  8.760 1.550 8.920 1.955 ;
        RECT  8.635 2.975 8.920 3.205 ;
        RECT  7.690 1.725 8.760 1.955 ;
        RECT  8.295 2.975 8.635 3.315 ;
        RECT  8.300 1.090 8.530 1.495 ;
        RECT  7.055 1.265 8.300 1.495 ;
        RECT  7.840 0.630 8.070 1.035 ;
        RECT  5.265 0.805 7.840 1.035 ;
        RECT  7.350 1.725 7.690 2.235 ;
        RECT  7.055 2.625 7.290 2.855 ;
        RECT  7.040 4.005 7.270 4.410 ;
        RECT  6.825 1.265 7.055 2.855 ;
        RECT  3.580 4.180 7.040 4.410 ;
        RECT  6.365 3.545 6.595 3.950 ;
        RECT  1.785 3.720 6.365 3.950 ;
        RECT  5.985 2.020 6.065 3.490 ;
        RECT  5.835 1.450 5.985 3.490 ;
        RECT  5.755 1.450 5.835 2.250 ;
        RECT  3.225 3.260 5.835 3.490 ;
        RECT  5.265 2.800 5.400 3.030 ;
        RECT  5.035 0.805 5.265 3.030 ;
        RECT  4.485 2.800 4.680 3.030 ;
        RECT  4.485 0.860 4.600 1.320 ;
        RECT  4.255 0.860 4.485 3.030 ;
        RECT  2.320 0.860 4.255 1.090 ;
        RECT  3.720 2.800 3.920 3.030 ;
        RECT  3.720 1.325 3.880 1.665 ;
        RECT  3.490 1.325 3.720 3.030 ;
        RECT  2.995 1.325 3.225 3.490 ;
        RECT  2.820 1.325 2.995 1.665 ;
        RECT  2.820 3.150 2.995 3.490 ;
        RECT  2.320 2.205 2.750 2.545 ;
        RECT  2.090 0.860 2.320 3.315 ;
        RECT  1.500 1.390 2.090 1.800 ;
        RECT  1.500 3.085 2.090 3.315 ;
        RECT  1.555 3.615 1.785 3.950 ;
        RECT  0.520 3.615 1.555 3.845 ;
        RECT  0.980 1.570 1.500 1.800 ;
        RECT  0.810 1.570 0.980 2.260 ;
        RECT  0.750 1.570 0.810 2.390 ;
        RECT  0.580 2.030 0.750 2.390 ;
        RECT  0.350 0.835 0.520 1.645 ;
        RECT  0.350 2.940 0.520 4.220 ;
        RECT  0.180 0.835 0.350 4.220 ;
        RECT  0.120 1.415 0.180 3.170 ;
    END
END AFCSHCINX4

MACRO AFCSHCINX2
    CLASS CORE ;
    FOREIGN AFCSHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFCSHCINX4 ;
    SIZE 33.000 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  32.715 2.940 32.860 4.340 ;
        RECT  32.715 0.970 32.770 1.845 ;
        RECT  32.485 0.970 32.715 4.340 ;
        RECT  32.480 0.970 32.485 1.820 ;
        RECT  32.480 2.940 32.485 4.340 ;
        RECT  32.430 0.970 32.480 1.780 ;
        RECT  32.380 2.940 32.480 4.220 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  31.655 1.260 32.200 1.540 ;
        RECT  31.425 1.260 31.655 2.465 ;
        RECT  31.235 2.120 31.425 2.465 ;
        RECT  31.180 2.120 31.235 2.460 ;
        END
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.775 3.425 22.040 3.765 ;
        RECT  21.775 1.475 21.885 1.815 ;
        RECT  21.640 1.475 21.775 3.765 ;
        RECT  21.545 1.475 21.640 3.780 ;
        RECT  21.260 2.940 21.545 3.780 ;
        RECT  20.990 3.425 21.260 3.780 ;
        RECT  20.760 3.425 20.990 3.875 ;
        RECT  19.860 3.645 20.760 3.875 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.430 3.260 18.220 3.490 ;
        RECT  16.430 1.690 16.540 1.920 ;
        RECT  16.200 1.690 16.430 3.490 ;
        RECT  15.950 2.940 16.200 3.490 ;
        RECT  15.945 2.940 15.950 3.365 ;
        END
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  25.700 2.300 26.260 2.780 ;
        END
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 2.055 9.915 2.660 ;
        END
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 2.245 8.685 2.700 ;
        RECT  7.860 2.470 8.060 2.700 ;
        RECT  7.630 2.470 7.860 3.315 ;
        RECT  6.595 3.085 7.630 3.315 ;
        RECT  6.515 2.035 6.595 3.440 ;
        RECT  6.365 1.390 6.515 3.440 ;
        RECT  6.285 1.390 6.365 2.265 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.490 2.105 1.600 2.445 ;
        RECT  1.260 2.105 1.490 2.850 ;
        RECT  1.180 2.620 1.260 2.850 ;
        RECT  0.950 2.620 1.180 3.195 ;
        RECT  0.875 2.965 0.950 3.195 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  32.010 -0.400 33.000 0.400 ;
        RECT  31.670 -0.400 32.010 0.630 ;
        RECT  30.435 -0.400 31.670 0.400 ;
        RECT  30.205 -0.400 30.435 1.760 ;
        RECT  27.370 -0.400 30.205 0.400 ;
        RECT  27.030 -0.400 27.370 0.575 ;
        RECT  25.195 -0.400 27.030 0.400 ;
        RECT  24.855 -0.400 25.195 0.575 ;
        RECT  13.060 -0.400 24.855 0.400 ;
        RECT  12.720 -0.400 13.060 0.575 ;
        RECT  6.695 -0.400 12.720 0.400 ;
        RECT  6.355 -0.400 6.695 0.575 ;
        RECT  2.400 -0.400 6.355 0.400 ;
        RECT  2.060 -0.400 2.400 0.575 ;
        RECT  1.280 -0.400 2.060 0.400 ;
        RECT  0.940 -0.400 1.280 0.630 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  31.960 4.640 33.000 5.440 ;
        RECT  31.620 3.760 31.960 5.440 ;
        RECT  31.160 4.640 31.620 5.440 ;
        RECT  30.820 3.760 31.160 5.440 ;
        RECT  27.360 4.640 30.820 5.440 ;
        RECT  27.020 3.150 27.360 5.440 ;
        RECT  25.430 4.640 27.020 5.440 ;
        RECT  25.090 4.465 25.430 5.440 ;
        RECT  10.960 4.640 25.090 5.440 ;
        RECT  10.620 4.465 10.960 5.440 ;
        RECT  9.395 4.640 10.620 5.440 ;
        RECT  9.055 4.465 9.395 5.440 ;
        RECT  8.090 4.640 9.055 5.440 ;
        RECT  7.750 4.465 8.090 5.440 ;
        RECT  2.390 4.640 7.750 5.440 ;
        RECT  2.050 4.465 2.390 5.440 ;
        RECT  1.240 4.640 2.050 5.440 ;
        RECT  0.900 4.080 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  32.115 2.170 32.225 2.510 ;
        RECT  31.885 2.170 32.115 3.530 ;
        RECT  30.590 3.300 31.885 3.530 ;
        RECT  30.950 2.840 31.200 3.070 ;
        RECT  30.950 1.460 31.190 1.800 ;
        RECT  30.720 1.460 30.950 3.070 ;
        RECT  30.130 2.840 30.720 3.070 ;
        RECT  30.360 3.300 30.590 4.405 ;
        RECT  28.745 4.175 30.360 4.405 ;
        RECT  29.900 2.840 30.130 3.915 ;
        RECT  29.745 0.805 29.975 2.355 ;
        RECT  29.205 3.685 29.900 3.915 ;
        RECT  20.255 0.805 29.745 1.035 ;
        RECT  29.515 2.670 29.670 3.450 ;
        RECT  29.440 1.380 29.515 3.450 ;
        RECT  29.285 1.380 29.440 2.900 ;
        RECT  29.000 3.130 29.205 3.915 ;
        RECT  28.975 2.170 29.000 3.915 ;
        RECT  28.770 2.170 28.975 3.360 ;
        RECT  28.540 1.380 28.850 1.720 ;
        RECT  28.540 3.595 28.745 4.405 ;
        RECT  28.515 1.380 28.540 4.405 ;
        RECT  28.310 1.380 28.515 3.825 ;
        RECT  28.075 3.110 28.080 4.390 ;
        RECT  27.845 1.460 28.075 4.390 ;
        RECT  27.740 3.110 27.845 4.390 ;
        RECT  27.440 2.270 27.550 2.610 ;
        RECT  27.210 1.270 27.440 2.610 ;
        RECT  23.660 1.270 27.210 1.500 ;
        RECT  26.490 1.730 26.720 4.410 ;
        RECT  26.270 1.730 26.490 1.960 ;
        RECT  26.260 3.710 26.490 4.410 ;
        RECT  23.200 3.710 26.260 3.940 ;
        RECT  25.455 3.020 25.990 3.250 ;
        RECT  25.455 1.730 25.910 1.960 ;
        RECT  25.225 1.730 25.455 3.250 ;
        RECT  24.620 2.260 25.225 2.490 ;
        RECT  24.560 3.140 24.670 3.480 ;
        RECT  24.380 2.780 24.560 3.480 ;
        RECT  24.380 1.730 24.440 1.960 ;
        RECT  24.330 1.730 24.380 3.480 ;
        RECT  24.150 1.730 24.330 3.010 ;
        RECT  22.545 4.180 24.320 4.410 ;
        RECT  24.095 1.730 24.150 1.960 ;
        RECT  23.660 3.250 23.950 3.480 ;
        RECT  23.430 1.270 23.660 3.480 ;
        RECT  22.970 1.670 23.200 3.940 ;
        RECT  22.605 1.670 22.970 1.900 ;
        RECT  22.890 3.710 22.970 3.940 ;
        RECT  22.545 2.240 22.740 2.825 ;
        RECT  22.265 1.560 22.605 1.900 ;
        RECT  22.510 2.240 22.545 4.410 ;
        RECT  22.315 2.595 22.510 4.410 ;
        RECT  11.420 4.180 22.315 4.410 ;
        RECT  21.055 1.415 21.165 1.755 ;
        RECT  20.825 1.415 21.055 2.435 ;
        RECT  19.865 2.205 20.825 2.435 ;
        RECT  20.025 0.805 20.255 1.885 ;
        RECT  19.405 1.655 20.025 1.885 ;
        RECT  19.635 2.205 19.865 3.415 ;
        RECT  18.365 1.080 19.645 1.420 ;
        RECT  19.490 3.185 19.635 3.415 ;
        RECT  19.140 3.185 19.490 3.950 ;
        RECT  19.175 1.655 19.405 2.955 ;
        RECT  17.000 2.725 19.175 2.955 ;
        RECT  11.880 3.720 19.140 3.950 ;
        RECT  17.460 2.265 18.940 2.495 ;
        RECT  17.230 0.770 17.460 2.495 ;
        RECT  13.825 0.770 17.230 1.000 ;
        RECT  16.770 1.230 17.000 2.955 ;
        RECT  15.250 1.230 16.770 1.460 ;
        RECT  15.710 1.690 15.820 1.920 ;
        RECT  15.480 1.690 15.710 3.490 ;
        RECT  12.340 3.260 15.480 3.490 ;
        RECT  15.020 1.230 15.250 3.030 ;
        RECT  14.720 1.230 15.020 1.570 ;
        RECT  14.090 2.800 15.020 3.030 ;
        RECT  14.055 1.230 14.285 2.565 ;
        RECT  13.860 2.335 14.055 2.565 ;
        RECT  13.630 2.335 13.860 3.030 ;
        RECT  13.595 0.770 13.825 1.565 ;
        RECT  13.370 2.800 13.630 3.030 ;
        RECT  12.030 1.335 13.595 1.565 ;
        RECT  12.490 0.875 13.210 1.105 ;
        RECT  12.910 2.120 13.190 2.350 ;
        RECT  12.570 2.120 12.910 3.030 ;
        RECT  11.570 2.120 12.570 2.350 ;
        RECT  12.260 0.630 12.490 1.105 ;
        RECT  12.110 3.085 12.340 3.490 ;
        RECT  7.155 0.630 12.260 0.860 ;
        RECT  10.430 3.085 12.110 3.315 ;
        RECT  11.800 1.090 12.030 1.565 ;
        RECT  11.650 3.545 11.880 3.950 ;
        RECT  7.615 1.090 11.800 1.320 ;
        RECT  7.055 3.545 11.650 3.775 ;
        RECT  11.340 1.550 11.570 2.350 ;
        RECT  11.190 4.005 11.420 4.410 ;
        RECT  11.230 1.550 11.340 1.780 ;
        RECT  7.520 4.005 11.190 4.235 ;
        RECT  10.200 1.550 10.430 3.315 ;
        RECT  9.970 1.550 10.200 1.780 ;
        RECT  9.815 2.975 10.200 3.315 ;
        RECT  8.920 1.550 9.150 3.205 ;
        RECT  8.080 1.550 8.920 1.780 ;
        RECT  8.635 2.975 8.920 3.205 ;
        RECT  8.295 2.975 8.635 3.315 ;
        RECT  7.850 1.550 8.080 1.955 ;
        RECT  7.830 1.725 7.850 1.955 ;
        RECT  7.490 1.725 7.830 2.165 ;
        RECT  7.385 1.090 7.615 1.495 ;
        RECT  7.290 4.005 7.520 4.410 ;
        RECT  7.260 1.265 7.385 1.495 ;
        RECT  3.580 4.180 7.290 4.410 ;
        RECT  7.030 1.265 7.260 2.855 ;
        RECT  6.925 0.630 7.155 1.035 ;
        RECT  6.825 3.545 7.055 3.950 ;
        RECT  6.825 2.625 7.030 2.855 ;
        RECT  5.265 0.805 6.925 1.035 ;
        RECT  1.710 3.720 6.825 3.950 ;
        RECT  5.985 2.495 6.065 3.490 ;
        RECT  5.835 1.265 5.985 3.490 ;
        RECT  5.755 1.265 5.835 2.725 ;
        RECT  3.225 3.260 5.835 3.490 ;
        RECT  5.265 2.800 5.400 3.030 ;
        RECT  5.035 0.805 5.265 3.030 ;
        RECT  4.485 2.800 4.680 3.030 ;
        RECT  4.485 0.860 4.600 1.320 ;
        RECT  4.255 0.860 4.485 3.030 ;
        RECT  2.320 0.860 4.255 1.090 ;
        RECT  3.720 2.800 3.920 3.030 ;
        RECT  3.720 1.325 3.880 1.665 ;
        RECT  3.490 1.325 3.720 3.030 ;
        RECT  2.995 1.325 3.225 3.490 ;
        RECT  2.820 1.325 2.995 1.665 ;
        RECT  2.820 3.150 2.995 3.490 ;
        RECT  2.320 2.205 2.750 2.545 ;
        RECT  2.090 0.860 2.320 3.315 ;
        RECT  1.500 1.390 2.090 1.800 ;
        RECT  1.500 3.085 2.090 3.315 ;
        RECT  1.480 3.590 1.710 3.950 ;
        RECT  0.980 1.570 1.500 1.800 ;
        RECT  0.520 3.590 1.480 3.820 ;
        RECT  0.810 1.570 0.980 2.260 ;
        RECT  0.750 1.570 0.810 2.390 ;
        RECT  0.580 2.030 0.750 2.390 ;
        RECT  0.350 0.835 0.520 1.645 ;
        RECT  0.350 2.940 0.520 4.220 ;
        RECT  0.180 0.835 0.350 4.220 ;
        RECT  0.120 1.415 0.180 3.170 ;
    END
END AFCSHCINX2

MACRO AHHCONX4
    CLASS CORE ;
    FOREIGN AHHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 1.820 4.480 3.220 ;
        RECT  4.100 1.330 4.330 3.220 ;
        RECT  3.935 1.330 4.100 1.560 ;
        RECT  3.515 2.840 4.100 3.070 ;
        RECT  3.615 1.210 3.935 1.560 ;
        RECT  3.500 2.840 3.515 3.220 ;
        RECT  3.270 2.840 3.500 3.685 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.420 1.820 8.440 3.220 ;
        RECT  8.060 1.365 8.420 3.430 ;
        RECT  6.815 1.365 8.060 1.595 ;
        RECT  7.445 3.090 8.060 3.430 ;
        RECT  7.105 3.090 7.445 3.900 ;
        RECT  5.960 3.090 7.105 3.430 ;
        RECT  6.700 1.260 6.815 1.595 ;
        RECT  6.360 0.705 6.700 1.595 ;
        RECT  5.640 3.090 5.960 3.900 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.095 2.290 6.940 2.690 ;
        RECT  5.410 2.460 6.095 2.690 ;
        RECT  5.180 2.460 5.410 4.145 ;
        RECT  3.040 3.915 5.180 4.145 ;
        RECT  3.640 1.800 3.870 2.520 ;
        RECT  3.040 2.290 3.640 2.520 ;
        RECT  2.810 2.290 3.040 4.145 ;
        RECT  2.215 2.290 2.810 2.660 ;
        RECT  1.875 2.235 2.215 2.660 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.345 1.830 7.685 2.230 ;
        RECT  5.725 1.830 7.345 2.060 ;
        RECT  5.660 1.285 5.725 2.060 ;
        RECT  5.495 1.285 5.660 2.230 ;
        RECT  5.320 1.830 5.495 2.230 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.020 -0.400 8.580 0.400 ;
        RECT  7.680 -0.400 8.020 1.105 ;
        RECT  5.380 -0.400 7.680 0.400 ;
        RECT  5.040 -0.400 5.380 0.575 ;
        RECT  1.340 -0.400 5.040 0.400 ;
        RECT  1.000 -0.400 1.340 0.575 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.245 4.640 8.580 5.440 ;
        RECT  7.905 3.935 8.245 5.440 ;
        RECT  6.685 4.640 7.905 5.440 ;
        RECT  6.345 3.935 6.685 5.440 ;
        RECT  5.035 4.640 6.345 5.440 ;
        RECT  4.695 4.410 5.035 5.440 ;
        RECT  1.335 4.640 4.695 5.440 ;
        RECT  0.995 4.410 1.335 5.440 ;
        RECT  0.000 4.640 0.995 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.720 0.810 4.950 3.685 ;
        RECT  4.620 0.810 4.720 1.040 ;
        RECT  3.935 3.455 4.720 3.685 ;
        RECT  4.280 0.675 4.620 1.040 ;
        RECT  3.385 0.730 4.280 0.960 ;
        RECT  3.155 0.730 3.385 1.955 ;
        RECT  1.490 1.725 3.155 1.955 ;
        RECT  2.600 0.630 2.925 1.035 ;
        RECT  1.030 1.265 2.680 1.495 ;
        RECT  0.570 0.805 2.600 1.035 ;
        RECT  2.215 3.920 2.530 4.290 ;
        RECT  0.570 3.920 2.215 4.150 ;
        RECT  1.705 3.180 2.045 3.520 ;
        RECT  1.030 3.180 1.705 3.410 ;
        RECT  1.260 1.725 1.490 2.560 ;
        RECT  0.800 1.265 1.030 3.410 ;
        RECT  0.230 0.760 0.570 4.150 ;
    END
END AHHCONX4

MACRO AHHCONX2
    CLASS CORE ;
    FOREIGN AHHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AHHCONX4 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.260 1.330 4.490 3.220 ;
        RECT  3.845 1.330 4.260 1.560 ;
        RECT  3.500 2.840 4.260 3.220 ;
        RECT  3.615 1.210 3.845 1.560 ;
        RECT  3.270 2.840 3.500 3.685 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.285 7.045 4.040 ;
        RECT  6.700 1.260 6.815 1.515 ;
        RECT  5.640 3.700 6.815 4.040 ;
        RECT  6.360 0.705 6.700 1.515 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.090 2.235 6.320 3.300 ;
        RECT  5.410 3.070 6.090 3.300 ;
        RECT  5.180 3.070 5.410 4.145 ;
        RECT  3.040 3.915 5.180 4.145 ;
        RECT  3.800 1.800 4.030 2.520 ;
        RECT  3.040 2.290 3.800 2.520 ;
        RECT  2.810 2.290 3.040 4.145 ;
        RECT  2.370 2.290 2.810 2.660 ;
        RECT  2.030 2.235 2.370 2.660 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.760 1.740 5.315 2.300 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 -0.400 7.260 0.400 ;
        RECT  5.040 -0.400 5.380 0.575 ;
        RECT  1.340 -0.400 5.040 0.400 ;
        RECT  1.000 -0.400 1.340 0.575 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.685 4.640 7.260 5.440 ;
        RECT  6.345 4.410 6.685 5.440 ;
        RECT  5.035 4.640 6.345 5.440 ;
        RECT  4.695 4.410 5.035 5.440 ;
        RECT  1.335 4.640 4.695 5.440 ;
        RECT  0.995 4.410 1.335 5.440 ;
        RECT  0.000 4.640 0.995 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.565 0.810 5.795 2.825 ;
        RECT  4.620 0.810 5.565 1.040 ;
        RECT  4.950 2.595 5.565 2.825 ;
        RECT  4.720 2.595 4.950 3.685 ;
        RECT  3.935 3.455 4.720 3.685 ;
        RECT  4.280 0.675 4.620 1.040 ;
        RECT  3.385 0.730 4.280 0.960 ;
        RECT  3.155 0.730 3.385 1.955 ;
        RECT  1.605 1.725 3.155 1.955 ;
        RECT  2.600 0.630 2.925 1.035 ;
        RECT  1.035 1.265 2.805 1.495 ;
        RECT  0.575 0.805 2.600 1.035 ;
        RECT  2.265 3.920 2.580 4.290 ;
        RECT  0.575 3.920 2.265 4.150 ;
        RECT  1.755 3.180 2.095 3.520 ;
        RECT  1.035 3.180 1.755 3.410 ;
        RECT  1.375 1.725 1.605 2.560 ;
        RECT  1.265 2.220 1.375 2.560 ;
        RECT  0.805 1.265 1.035 3.410 ;
        RECT  0.235 0.760 0.575 4.150 ;
    END
END AHHCONX2

MACRO AHHCINX4
    CLASS CORE ;
    FOREIGN AHHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.215 2.910 3.555 3.730 ;
        RECT  3.180 1.270 3.410 2.050 ;
        RECT  3.160 2.910 3.215 3.220 ;
        RECT  3.160 1.820 3.180 2.050 ;
        RECT  2.780 1.820 3.160 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.320 1.260 8.440 2.780 ;
        RECT  8.060 0.990 8.320 2.780 ;
        RECT  7.980 0.990 8.060 1.800 ;
        RECT  7.720 2.550 8.060 2.780 ;
        RECT  7.780 1.260 7.980 1.560 ;
        RECT  6.925 1.330 7.780 1.560 ;
        RECT  7.380 2.550 7.720 3.590 ;
        RECT  6.585 0.730 6.925 1.560 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.900 2.130 9.010 2.470 ;
        RECT  8.670 2.130 8.900 3.240 ;
        RECT  8.180 3.010 8.670 3.240 ;
        RECT  7.950 3.010 8.180 4.130 ;
        RECT  6.625 3.900 7.950 4.130 ;
        RECT  6.395 2.250 6.625 4.130 ;
        RECT  4.405 3.900 6.395 4.130 ;
        RECT  4.175 3.900 4.405 4.370 ;
        RECT  1.510 4.140 4.175 4.370 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.140 1.990 5.165 2.330 ;
        RECT  4.760 1.990 5.140 2.660 ;
        RECT  4.355 1.990 4.760 2.330 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 -0.400 9.240 0.400 ;
        RECT  8.700 -0.400 9.040 1.800 ;
        RECT  7.685 -0.400 8.700 0.400 ;
        RECT  7.345 -0.400 7.685 0.630 ;
        RECT  6.165 -0.400 7.345 0.400 ;
        RECT  5.825 -0.400 6.165 0.575 ;
        RECT  4.905 -0.400 5.825 0.400 ;
        RECT  4.565 -0.400 4.905 1.250 ;
        RECT  1.280 -0.400 4.565 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 4.640 9.240 5.440 ;
        RECT  8.700 3.470 9.040 5.440 ;
        RECT  6.350 4.640 8.700 5.440 ;
        RECT  6.010 4.465 6.350 5.440 ;
        RECT  5.080 4.640 6.010 5.440 ;
        RECT  4.740 4.465 5.080 5.440 ;
        RECT  1.280 4.640 4.740 5.440 ;
        RECT  0.940 4.410 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.200 2.045 7.820 2.275 ;
        RECT  6.970 1.790 7.200 2.275 ;
        RECT  5.740 1.790 6.970 2.020 ;
        RECT  5.740 2.760 5.795 3.580 ;
        RECT  5.625 1.790 5.740 3.580 ;
        RECT  5.510 1.270 5.625 3.580 ;
        RECT  5.395 1.270 5.510 2.020 ;
        RECT  5.455 2.760 5.510 3.580 ;
        RECT  5.285 1.270 5.395 1.610 ;
        RECT  4.125 2.910 4.285 3.670 ;
        RECT  4.125 0.765 4.185 1.575 ;
        RECT  3.895 0.765 4.125 3.670 ;
        RECT  3.845 0.765 3.895 1.575 ;
        RECT  2.950 0.765 3.845 0.995 ;
        RECT  2.720 0.765 2.950 1.495 ;
        RECT  2.455 3.570 2.795 3.910 ;
        RECT  2.405 1.265 2.720 1.495 ;
        RECT  2.180 0.630 2.490 1.035 ;
        RECT  0.520 3.680 2.455 3.910 ;
        RECT  2.085 2.230 2.425 2.570 ;
        RECT  2.175 1.265 2.405 1.955 ;
        RECT  0.520 0.805 2.180 1.035 ;
        RECT  1.270 1.725 2.175 1.955 ;
        RECT  1.880 2.340 2.085 2.570 ;
        RECT  1.650 2.340 1.880 3.450 ;
        RECT  0.810 1.265 1.845 1.495 ;
        RECT  1.540 2.800 1.650 3.450 ;
        RECT  0.810 2.800 1.540 3.030 ;
        RECT  1.040 1.725 1.270 2.500 ;
        RECT  0.580 1.265 0.810 3.030 ;
        RECT  0.350 0.695 0.520 1.035 ;
        RECT  0.350 3.375 0.520 4.185 ;
        RECT  0.120 0.695 0.350 4.185 ;
    END
END AHHCINX4

MACRO AHHCINX2
    CLASS CORE ;
    FOREIGN AHHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AHHCINX4 ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.215 2.910 3.555 3.730 ;
        RECT  3.180 1.210 3.410 1.955 ;
        RECT  3.095 2.910 3.215 3.220 ;
        RECT  3.095 1.725 3.180 1.955 ;
        RECT  2.865 1.725 3.095 3.220 ;
        RECT  2.855 2.405 2.865 2.635 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.675 2.405 7.705 3.755 ;
        RECT  7.525 1.330 7.675 3.755 ;
        RECT  7.445 1.330 7.525 4.060 ;
        RECT  6.855 1.330 7.445 1.560 ;
        RECT  7.355 2.380 7.445 4.060 ;
        RECT  7.185 2.780 7.355 4.060 ;
        RECT  6.515 0.630 6.855 1.560 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.170 2.250 6.400 3.710 ;
        RECT  4.410 3.480 6.170 3.710 ;
        RECT  4.180 3.480 4.410 4.370 ;
        RECT  4.175 4.085 4.180 4.370 ;
        RECT  1.510 4.140 4.175 4.370 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.065 1.800 5.080 2.140 ;
        RECT  4.835 1.800 5.065 2.635 ;
        RECT  4.740 1.800 4.835 2.140 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.615 -0.400 7.920 0.400 ;
        RECT  7.275 -0.400 7.615 1.100 ;
        RECT  6.095 -0.400 7.275 0.400 ;
        RECT  5.755 -0.400 6.095 0.575 ;
        RECT  4.945 -0.400 5.755 0.400 ;
        RECT  4.605 -0.400 4.945 0.575 ;
        RECT  1.285 -0.400 4.605 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.180 4.640 7.920 5.440 ;
        RECT  5.840 3.940 6.180 5.440 ;
        RECT  5.050 4.640 5.840 5.440 ;
        RECT  4.710 3.940 5.050 5.440 ;
        RECT  1.280 4.640 4.710 5.440 ;
        RECT  0.940 4.410 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.815 1.790 7.155 2.130 ;
        RECT  5.600 1.790 6.815 2.020 ;
        RECT  5.370 1.170 5.600 3.250 ;
        RECT  5.205 1.170 5.370 1.510 ;
        RECT  5.255 2.910 5.370 3.250 ;
        RECT  4.220 2.910 4.275 3.250 ;
        RECT  3.990 0.700 4.220 3.250 ;
        RECT  3.845 0.700 3.990 1.510 ;
        RECT  3.935 2.910 3.990 3.250 ;
        RECT  2.950 0.700 3.845 0.930 ;
        RECT  2.720 0.700 2.950 1.495 ;
        RECT  2.405 1.265 2.720 1.495 ;
        RECT  2.295 3.100 2.635 3.910 ;
        RECT  2.165 0.630 2.490 1.035 ;
        RECT  2.085 2.230 2.425 2.570 ;
        RECT  2.175 1.265 2.405 1.955 ;
        RECT  0.520 3.680 2.295 3.910 ;
        RECT  1.270 1.725 2.175 1.955 ;
        RECT  0.520 0.805 2.165 1.035 ;
        RECT  1.880 2.340 2.085 2.570 ;
        RECT  1.650 2.340 1.880 3.450 ;
        RECT  0.810 1.265 1.845 1.495 ;
        RECT  1.540 2.770 1.650 3.450 ;
        RECT  0.810 2.770 1.540 3.000 ;
        RECT  1.040 1.725 1.270 2.500 ;
        RECT  0.580 1.265 0.810 3.000 ;
        RECT  0.350 0.695 0.520 1.035 ;
        RECT  0.350 3.375 0.520 4.185 ;
        RECT  0.120 0.695 0.350 4.185 ;
    END
END AHHCINX2

MACRO AFHCONX4
    CLASS CORE ;
    FOREIGN AFHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.000 2.940 17.020 4.340 ;
        RECT  16.975 2.635 17.000 4.340 ;
        RECT  16.975 0.940 16.980 1.875 ;
        RECT  16.640 0.940 16.975 4.340 ;
        RECT  16.635 1.200 16.640 3.040 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.330 0.680 10.670 1.020 ;
        RECT  9.300 0.790 10.330 1.020 ;
        RECT  9.760 2.800 9.965 3.030 ;
        RECT  9.610 1.820 9.760 3.220 ;
        RECT  9.380 1.820 9.610 3.480 ;
        RECT  9.300 1.820 9.380 2.050 ;
        RECT  8.675 3.250 9.380 3.480 ;
        RECT  9.070 0.790 9.300 2.050 ;
        RECT  8.505 1.270 9.070 1.610 ;
        RECT  8.445 3.250 8.675 4.350 ;
        RECT  8.185 4.010 8.445 4.350 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.400 2.000 14.210 2.640 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 2.135 7.145 2.790 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.215 0.830 2.635 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.190 -0.400 17.160 0.400 ;
        RECT  15.850 -0.400 16.190 0.575 ;
        RECT  14.830 -0.400 15.850 0.400 ;
        RECT  14.490 -0.400 14.830 0.575 ;
        RECT  13.470 -0.400 14.490 0.400 ;
        RECT  13.130 -0.400 13.470 0.575 ;
        RECT  7.000 -0.400 13.130 0.400 ;
        RECT  6.660 -0.400 7.000 0.575 ;
        RECT  1.285 -0.400 6.660 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.915 4.640 17.160 5.440 ;
        RECT  15.575 3.940 15.915 5.440 ;
        RECT  14.505 4.640 15.575 5.440 ;
        RECT  14.165 4.465 14.505 5.440 ;
        RECT  13.145 4.640 14.165 5.440 ;
        RECT  12.805 4.465 13.145 5.440 ;
        RECT  7.020 4.640 12.805 5.440 ;
        RECT  6.680 4.090 7.020 5.440 ;
        RECT  1.325 4.640 6.680 5.440 ;
        RECT  0.985 3.620 1.325 5.440 ;
        RECT  0.000 4.640 0.985 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.340 2.040 16.365 2.550 ;
        RECT  16.135 0.895 16.340 2.550 ;
        RECT  16.110 0.895 16.135 2.270 ;
        RECT  14.675 0.895 16.110 1.125 ;
        RECT  15.400 1.360 15.510 1.700 ;
        RECT  15.170 1.360 15.400 2.320 ;
        RECT  15.135 2.090 15.170 2.320 ;
        RECT  14.905 2.090 15.135 4.215 ;
        RECT  11.550 3.985 14.905 4.215 ;
        RECT  14.445 0.895 14.675 3.740 ;
        RECT  11.570 3.510 14.445 3.740 ;
        RECT  13.810 1.360 14.150 1.700 ;
        RECT  13.485 2.930 13.825 3.270 ;
        RECT  13.170 1.415 13.810 1.645 ;
        RECT  13.105 2.985 13.485 3.215 ;
        RECT  13.105 0.825 13.170 2.100 ;
        RECT  12.940 0.825 13.105 3.215 ;
        RECT  12.490 0.825 12.940 1.055 ;
        RECT  12.875 1.865 12.940 3.215 ;
        RECT  12.575 2.230 12.875 2.460 ;
        RECT  12.450 1.340 12.710 1.570 ;
        RECT  12.260 0.630 12.490 1.055 ;
        RECT  12.280 1.340 12.450 1.945 ;
        RECT  12.280 2.805 12.335 3.145 ;
        RECT  12.220 1.340 12.280 3.145 ;
        RECT  11.270 0.630 12.260 0.860 ;
        RECT  12.050 1.715 12.220 3.145 ;
        RECT  11.995 2.805 12.050 3.145 ;
        RECT  11.755 1.095 11.990 1.435 ;
        RECT  11.570 1.095 11.755 2.515 ;
        RECT  11.525 1.095 11.570 3.740 ;
        RECT  11.320 3.985 11.550 4.410 ;
        RECT  11.340 2.285 11.525 3.740 ;
        RECT  11.230 2.850 11.340 3.740 ;
        RECT  10.230 4.180 11.320 4.410 ;
        RECT  11.040 0.630 11.270 1.800 ;
        RECT  10.985 1.460 11.040 1.800 ;
        RECT  10.755 1.460 10.985 3.950 ;
        RECT  10.470 3.720 10.755 3.950 ;
        RECT  10.230 1.300 10.440 3.490 ;
        RECT  10.210 1.300 10.230 4.410 ;
        RECT  9.610 1.300 10.210 1.530 ;
        RECT  10.000 3.260 10.210 4.410 ;
        RECT  9.245 3.895 10.000 4.130 ;
        RECT  8.905 3.790 9.245 4.130 ;
        RECT  8.605 2.205 8.835 3.020 ;
        RECT  8.570 0.645 8.800 1.035 ;
        RECT  8.215 2.790 8.605 3.020 ;
        RECT  8.245 0.805 8.570 1.035 ;
        RECT  8.015 0.805 8.245 2.560 ;
        RECT  7.985 2.790 8.215 3.780 ;
        RECT  6.205 0.805 8.015 1.035 ;
        RECT  7.880 2.220 8.015 2.560 ;
        RECT  5.530 3.550 7.985 3.780 ;
        RECT  7.630 1.265 7.765 1.495 ;
        RECT  7.630 2.980 7.740 3.320 ;
        RECT  7.400 1.265 7.630 3.320 ;
        RECT  6.125 2.980 6.295 3.320 ;
        RECT  6.125 1.320 6.235 1.660 ;
        RECT  5.975 0.630 6.205 1.035 ;
        RECT  5.895 1.320 6.125 3.320 ;
        RECT  4.150 0.630 5.975 0.860 ;
        RECT  5.760 2.180 5.895 2.545 ;
        RECT  5.300 1.090 5.530 3.780 ;
        RECT  4.610 1.090 5.300 1.320 ;
        RECT  4.840 1.550 5.070 4.350 ;
        RECT  2.045 4.120 4.840 4.350 ;
        RECT  4.380 1.090 4.610 3.775 ;
        RECT  2.765 3.545 4.380 3.775 ;
        RECT  3.920 0.630 4.150 3.305 ;
        RECT  3.375 0.900 3.485 1.415 ;
        RECT  3.375 2.970 3.485 3.310 ;
        RECT  3.145 0.900 3.375 3.310 ;
        RECT  1.315 0.900 3.145 1.130 ;
        RECT  2.710 1.390 2.765 1.730 ;
        RECT  2.710 3.435 2.765 3.775 ;
        RECT  2.480 1.390 2.710 3.775 ;
        RECT  2.425 1.390 2.480 1.730 ;
        RECT  2.425 3.435 2.480 3.775 ;
        RECT  1.990 1.390 2.045 1.730 ;
        RECT  1.990 3.455 2.045 4.350 ;
        RECT  1.760 1.390 1.990 4.350 ;
        RECT  1.705 1.390 1.760 1.730 ;
        RECT  1.705 3.455 1.760 4.350 ;
        RECT  1.315 2.040 1.465 2.405 ;
        RECT  1.085 0.900 1.315 3.180 ;
        RECT  0.525 1.345 1.085 1.575 ;
        RECT  0.605 2.950 1.085 3.180 ;
        RECT  0.265 2.950 0.605 4.230 ;
        RECT  0.185 0.765 0.525 1.575 ;
    END
END AFHCONX4

MACRO AFHCONX2
    CLASS CORE ;
    FOREIGN AFHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFHCONX4 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.370 0.965 13.480 1.775 ;
        RECT  13.140 0.965 13.370 3.020 ;
        RECT  13.115 2.790 13.140 3.020 ;
        RECT  12.870 2.790 13.115 3.250 ;
        RECT  12.755 2.790 12.870 3.195 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.945 1.215 9.175 3.535 ;
        RECT  8.330 1.215 8.945 1.555 ;
        RECT  8.560 3.305 8.945 3.535 ;
        RECT  8.330 3.305 8.560 4.225 ;
        RECT  8.020 3.995 8.330 4.225 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.965 1.940 15.075 2.570 ;
        RECT  14.675 1.845 14.965 2.570 ;
        RECT  14.435 1.940 14.675 2.570 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.340 2.140 7.120 2.695 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.215 2.110 0.760 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.900 -0.400 15.840 0.400 ;
        RECT  14.560 -0.400 14.900 1.590 ;
        RECT  12.720 -0.400 14.560 0.400 ;
        RECT  12.380 -0.400 12.720 0.575 ;
        RECT  6.880 -0.400 12.380 0.400 ;
        RECT  6.540 -0.400 6.880 0.575 ;
        RECT  1.280 -0.400 6.540 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.900 4.640 15.840 5.440 ;
        RECT  14.560 4.465 14.900 5.440 ;
        RECT  12.355 4.640 14.560 5.440 ;
        RECT  12.015 4.465 12.355 5.440 ;
        RECT  6.920 4.640 12.015 5.440 ;
        RECT  6.580 4.090 6.920 5.440 ;
        RECT  1.240 4.640 6.580 5.440 ;
        RECT  0.900 3.620 1.240 5.440 ;
        RECT  0.000 4.640 0.900 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.605 2.950 15.660 4.230 ;
        RECT  15.605 0.835 15.625 1.645 ;
        RECT  15.375 0.835 15.605 4.230 ;
        RECT  15.285 0.835 15.375 1.645 ;
        RECT  15.320 2.950 15.375 4.230 ;
        RECT  9.635 4.000 15.320 4.230 ;
        RECT  14.125 0.845 14.180 1.655 ;
        RECT  14.125 2.900 14.140 3.710 ;
        RECT  13.895 0.845 14.125 3.710 ;
        RECT  13.840 0.845 13.895 1.655 ;
        RECT  13.800 2.900 13.895 3.710 ;
        RECT  12.145 3.480 13.800 3.710 ;
        RECT  12.820 1.990 12.875 2.330 ;
        RECT  12.590 0.805 12.820 2.330 ;
        RECT  11.240 0.805 12.590 1.035 ;
        RECT  12.535 1.990 12.590 2.330 ;
        RECT  12.145 2.200 12.200 2.540 ;
        RECT  11.915 2.200 12.145 3.710 ;
        RECT  11.810 1.265 11.960 1.495 ;
        RECT  11.860 2.200 11.915 2.540 ;
        RECT  10.095 3.480 11.915 3.710 ;
        RECT  11.590 1.265 11.810 1.970 ;
        RECT  11.580 1.265 11.590 3.215 ;
        RECT  11.360 1.740 11.580 3.215 ;
        RECT  11.250 2.875 11.360 3.215 ;
        RECT  11.110 0.805 11.240 1.510 ;
        RECT  11.010 0.805 11.110 2.520 ;
        RECT  10.880 1.170 11.010 2.520 ;
        RECT  10.870 2.290 10.880 2.520 ;
        RECT  10.640 2.290 10.870 3.220 ;
        RECT  10.530 2.880 10.640 3.220 ;
        RECT  10.180 1.000 10.520 1.810 ;
        RECT  10.095 1.580 10.180 1.810 ;
        RECT  9.865 1.580 10.095 3.710 ;
        RECT  9.635 1.010 9.820 1.350 ;
        RECT  9.405 1.010 9.635 4.230 ;
        RECT  9.130 3.945 9.405 4.230 ;
        RECT  8.790 3.945 9.130 4.285 ;
        RECT  8.045 0.630 8.730 0.860 ;
        RECT  8.485 2.210 8.715 3.075 ;
        RECT  8.100 2.845 8.485 3.075 ;
        RECT  7.870 2.845 8.100 3.765 ;
        RECT  7.815 0.630 8.045 2.570 ;
        RECT  5.445 3.535 7.870 3.765 ;
        RECT  6.175 0.805 7.815 1.035 ;
        RECT  7.585 2.960 7.640 3.300 ;
        RECT  7.355 1.265 7.585 3.300 ;
        RECT  7.300 2.960 7.355 3.300 ;
        RECT  6.010 2.890 6.200 3.230 ;
        RECT  5.945 0.630 6.175 1.035 ;
        RECT  6.010 1.410 6.120 1.750 ;
        RECT  5.780 1.410 6.010 3.230 ;
        RECT  4.065 0.630 5.945 0.860 ;
        RECT  5.675 2.360 5.780 2.745 ;
        RECT  5.215 1.090 5.445 3.765 ;
        RECT  4.525 1.090 5.215 1.320 ;
        RECT  4.755 1.550 4.985 4.410 ;
        RECT  1.960 4.180 4.755 4.410 ;
        RECT  4.295 1.090 4.525 3.950 ;
        RECT  2.705 3.720 4.295 3.950 ;
        RECT  3.835 0.630 4.065 3.360 ;
        RECT  3.345 1.075 3.480 1.415 ;
        RECT  3.345 3.020 3.400 3.360 ;
        RECT  3.115 0.865 3.345 3.360 ;
        RECT  0.520 0.865 3.115 1.095 ;
        RECT  3.060 3.020 3.115 3.360 ;
        RECT  2.705 1.390 2.760 1.730 ;
        RECT  2.475 1.390 2.705 3.950 ;
        RECT  2.420 1.390 2.475 1.730 ;
        RECT  2.340 3.425 2.475 3.765 ;
        RECT  1.960 1.390 2.040 1.730 ;
        RECT  1.730 1.390 1.960 4.410 ;
        RECT  1.700 1.390 1.730 1.730 ;
        RECT  1.620 3.405 1.730 4.410 ;
        RECT  1.145 1.510 1.375 3.180 ;
        RECT  0.520 1.510 1.145 1.740 ;
        RECT  0.520 2.950 1.145 3.180 ;
        RECT  0.180 0.865 0.520 1.740 ;
        RECT  0.180 2.950 0.520 4.230 ;
    END
END AFHCONX2

MACRO AFHCINX4
    CLASS CORE ;
    FOREIGN AFHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.130 0.730 18.360 4.340 ;
        RECT  17.860 0.730 18.130 1.540 ;
        RECT  17.960 2.940 18.130 4.340 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.650 1.090 10.110 1.320 ;
        RECT  9.760 2.845 9.875 3.760 ;
        RECT  9.380 2.380 9.760 3.780 ;
        RECT  8.795 3.530 9.380 3.760 ;
        RECT  8.650 3.500 8.795 3.760 ;
        RECT  8.485 1.090 8.650 3.760 ;
        RECT  8.420 1.090 8.485 3.850 ;
        RECT  8.325 1.090 8.420 1.465 ;
        RECT  8.365 2.965 8.420 3.850 ;
        RECT  8.145 3.040 8.365 3.850 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 2.260 13.175 2.490 ;
        RECT  12.020 2.260 12.400 2.660 ;
        RECT  11.400 2.260 12.020 2.490 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.410 4.060 6.310 4.405 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.170 0.615 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.440 -0.400 18.480 0.400 ;
        RECT  17.100 -0.400 17.440 0.575 ;
        RECT  14.410 -0.400 17.100 0.400 ;
        RECT  14.070 -0.400 14.410 0.575 ;
        RECT  12.890 -0.400 14.070 0.400 ;
        RECT  12.550 -0.400 12.890 0.575 ;
        RECT  11.370 -0.400 12.550 0.400 ;
        RECT  11.030 -0.400 11.370 0.575 ;
        RECT  6.915 -0.400 11.030 0.400 ;
        RECT  6.575 -0.400 6.915 0.575 ;
        RECT  1.285 -0.400 6.575 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.335 4.640 18.480 5.440 ;
        RECT  16.525 4.465 17.335 5.440 ;
        RECT  13.780 4.640 16.525 5.440 ;
        RECT  13.420 4.395 13.780 5.440 ;
        RECT  12.285 4.640 13.420 5.440 ;
        RECT  11.945 3.860 12.285 5.440 ;
        RECT  10.805 4.640 11.945 5.440 ;
        RECT  10.465 4.465 10.805 5.440 ;
        RECT  7.040 4.640 10.465 5.440 ;
        RECT  6.700 4.090 7.040 5.440 ;
        RECT  1.325 4.640 6.700 5.440 ;
        RECT  0.985 3.610 1.325 5.440 ;
        RECT  0.000 4.640 0.985 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.730 2.035 17.900 2.710 ;
        RECT  17.670 2.035 17.730 4.170 ;
        RECT  17.500 2.480 17.670 4.170 ;
        RECT  15.530 3.940 17.500 4.170 ;
        RECT  17.000 0.835 17.230 2.250 ;
        RECT  15.320 0.835 17.000 1.065 ;
        RECT  16.540 1.295 16.770 3.600 ;
        RECT  16.335 1.295 16.540 1.635 ;
        RECT  16.100 3.370 16.540 3.600 ;
        RECT  16.080 1.865 16.310 3.140 ;
        RECT  15.760 3.370 16.100 3.710 ;
        RECT  15.940 1.865 16.080 2.095 ;
        RECT  15.530 2.910 16.080 3.140 ;
        RECT  15.710 1.295 15.940 2.095 ;
        RECT  15.620 2.325 15.850 2.680 ;
        RECT  15.600 1.295 15.710 1.635 ;
        RECT  14.740 2.325 15.620 2.555 ;
        RECT  15.300 2.910 15.530 4.170 ;
        RECT  15.090 0.835 15.320 1.675 ;
        RECT  14.655 3.645 15.300 3.985 ;
        RECT  13.795 1.445 15.090 1.675 ;
        RECT  14.150 0.895 14.840 1.125 ;
        RECT  14.510 2.060 14.740 3.415 ;
        RECT  14.380 2.060 14.510 2.400 ;
        RECT  13.725 3.185 14.510 3.415 ;
        RECT  13.795 2.725 14.275 2.955 ;
        RECT  13.920 0.805 14.150 1.125 ;
        RECT  10.630 0.805 13.920 1.035 ;
        RECT  13.650 1.445 13.795 2.955 ;
        RECT  13.495 3.185 13.725 3.630 ;
        RECT  13.565 1.390 13.650 2.955 ;
        RECT  13.310 1.390 13.565 1.730 ;
        RECT  13.005 2.725 13.565 2.955 ;
        RECT  10.335 3.400 13.495 3.630 ;
        RECT  12.775 2.725 13.005 3.170 ;
        RECT  12.665 2.830 12.775 3.170 ;
        RECT  11.790 1.385 12.130 1.780 ;
        RECT  11.155 1.550 11.790 1.780 ;
        RECT  11.225 2.830 11.565 3.170 ;
        RECT  11.155 2.830 11.225 3.060 ;
        RECT  10.925 1.550 11.155 3.060 ;
        RECT  10.830 1.550 10.925 1.780 ;
        RECT  10.490 1.390 10.830 1.780 ;
        RECT  10.400 0.630 10.630 1.035 ;
        RECT  9.150 1.550 10.490 1.780 ;
        RECT  8.095 0.630 10.400 0.860 ;
        RECT  10.235 2.310 10.335 4.220 ;
        RECT  10.105 2.310 10.235 4.310 ;
        RECT  10.005 3.990 10.105 4.310 ;
        RECT  7.605 4.080 10.005 4.310 ;
        RECT  8.920 1.550 9.150 3.265 ;
        RECT  7.865 0.630 8.095 2.585 ;
        RECT  6.140 0.805 7.865 1.035 ;
        RECT  7.635 3.025 7.765 3.365 ;
        RECT  7.405 1.275 7.635 3.365 ;
        RECT  7.375 3.595 7.605 4.310 ;
        RECT  5.610 3.595 7.375 3.825 ;
        RECT  6.945 2.165 7.175 2.530 ;
        RECT  6.100 2.165 6.945 2.395 ;
        RECT  6.075 2.980 6.320 3.320 ;
        RECT  5.910 0.630 6.140 1.035 ;
        RECT  6.075 1.335 6.100 2.395 ;
        RECT  5.870 1.335 6.075 3.320 ;
        RECT  4.230 0.630 5.910 0.860 ;
        RECT  5.845 2.165 5.870 3.320 ;
        RECT  5.380 1.090 5.610 3.825 ;
        RECT  4.690 1.090 5.380 1.320 ;
        RECT  4.920 1.550 5.150 4.335 ;
        RECT  2.045 4.105 4.920 4.335 ;
        RECT  4.460 1.090 4.690 3.795 ;
        RECT  2.805 3.565 4.460 3.795 ;
        RECT  4.000 0.630 4.230 3.300 ;
        RECT  3.225 0.930 3.565 3.300 ;
        RECT  1.245 0.930 3.225 1.160 ;
        RECT  2.465 1.390 2.805 3.795 ;
        RECT  2.460 2.990 2.465 3.795 ;
        RECT  1.815 1.390 2.045 4.335 ;
        RECT  1.705 1.390 1.815 1.730 ;
        RECT  1.705 3.405 1.815 4.335 ;
        RECT  1.245 2.015 1.580 2.405 ;
        RECT  1.015 0.930 1.245 3.170 ;
        RECT  0.525 1.475 1.015 1.705 ;
        RECT  0.605 2.940 1.015 3.170 ;
        RECT  0.265 2.940 0.605 4.220 ;
        RECT  0.185 0.765 0.525 1.705 ;
    END
END AFHCINX4

MACRO AFHCINX2
    CLASS CORE ;
    FOREIGN AFHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFHCINX4 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.285 2.940 16.360 4.340 ;
        RECT  16.140 1.335 16.285 4.340 ;
        RECT  16.055 0.730 16.140 4.340 ;
        RECT  15.800 0.730 16.055 1.565 ;
        RECT  15.980 2.940 16.055 4.340 ;
        RECT  15.685 3.110 15.980 3.920 ;
        RECT  15.795 1.020 15.800 1.565 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.885 1.110 10.120 1.450 ;
        RECT  9.655 1.110 9.885 1.980 ;
        RECT  9.450 1.750 9.655 1.980 ;
        RECT  9.320 1.750 9.450 3.755 ;
        RECT  9.220 1.750 9.320 3.780 ;
        RECT  8.720 3.500 9.220 3.780 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.675 2.195 11.430 2.660 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.620 2.940 7.780 3.220 ;
        RECT  7.615 2.220 7.620 3.220 ;
        RECT  7.385 2.220 7.615 3.760 ;
        RECT  7.175 2.220 7.385 2.560 ;
        RECT  6.130 3.530 7.385 3.760 ;
        RECT  5.900 1.095 6.130 3.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 2.170 0.615 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.380 -0.400 16.500 0.400 ;
        RECT  15.040 -0.400 15.380 0.575 ;
        RECT  11.635 -0.400 15.040 0.400 ;
        RECT  11.295 -0.400 11.635 0.575 ;
        RECT  7.665 -0.400 11.295 0.400 ;
        RECT  7.325 -0.400 7.665 0.575 ;
        RECT  1.285 -0.400 7.325 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.785 4.640 16.500 5.440 ;
        RECT  14.445 4.465 14.785 5.440 ;
        RECT  11.185 4.640 14.445 5.440 ;
        RECT  10.845 4.465 11.185 5.440 ;
        RECT  7.940 4.640 10.845 5.440 ;
        RECT  7.600 4.465 7.940 5.440 ;
        RECT  1.325 4.640 7.600 5.440 ;
        RECT  0.985 3.610 1.325 5.440 ;
        RECT  0.000 4.640 0.985 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.560 2.035 15.790 2.660 ;
        RECT  15.115 2.430 15.560 2.660 ;
        RECT  14.890 0.835 15.120 2.200 ;
        RECT  14.885 2.430 15.115 4.105 ;
        RECT  14.605 0.835 14.890 1.065 ;
        RECT  13.020 3.875 14.885 4.105 ;
        RECT  14.425 1.295 14.655 3.645 ;
        RECT  14.375 0.640 14.605 1.065 ;
        RECT  14.275 1.295 14.425 1.635 ;
        RECT  13.445 3.415 14.425 3.645 ;
        RECT  13.260 0.640 14.375 0.870 ;
        RECT  13.965 1.875 14.195 3.185 ;
        RECT  13.880 1.875 13.965 2.105 ;
        RECT  13.020 2.955 13.965 3.185 ;
        RECT  13.650 1.200 13.880 2.105 ;
        RECT  13.505 2.340 13.735 2.725 ;
        RECT  13.540 1.200 13.650 1.540 ;
        RECT  12.370 2.495 13.505 2.725 ;
        RECT  13.030 0.640 13.260 1.495 ;
        RECT  11.890 1.265 13.030 1.495 ;
        RECT  12.790 2.955 13.020 4.105 ;
        RECT  12.585 3.695 12.790 4.105 ;
        RECT  12.630 0.630 12.780 0.860 ;
        RECT  12.400 0.630 12.630 1.035 ;
        RECT  10.840 0.805 12.400 1.035 ;
        RECT  12.355 2.495 12.370 2.910 ;
        RECT  12.125 2.495 12.355 4.225 ;
        RECT  9.910 3.995 12.125 4.225 ;
        RECT  11.660 1.265 11.890 3.520 ;
        RECT  10.610 0.640 10.840 1.035 ;
        RECT  10.730 1.315 10.840 1.655 ;
        RECT  10.500 1.315 10.730 1.945 ;
        RECT  8.130 0.640 10.610 0.870 ;
        RECT  10.370 1.715 10.500 1.945 ;
        RECT  10.140 1.715 10.370 3.755 ;
        RECT  9.680 2.210 9.910 4.315 ;
        RECT  8.430 4.085 9.680 4.315 ;
        RECT  8.730 1.255 9.400 1.485 ;
        RECT  8.730 2.845 8.785 3.185 ;
        RECT  8.500 1.255 8.730 3.185 ;
        RECT  8.220 1.285 8.500 1.515 ;
        RECT  8.445 2.845 8.500 3.185 ;
        RECT  8.200 3.995 8.430 4.315 ;
        RECT  8.115 2.190 8.225 2.530 ;
        RECT  5.670 3.995 8.200 4.225 ;
        RECT  7.900 0.640 8.130 1.035 ;
        RECT  7.885 1.745 8.115 2.530 ;
        RECT  6.890 0.805 7.900 1.035 ;
        RECT  6.905 1.745 7.885 1.975 ;
        RECT  6.795 2.905 7.070 3.245 ;
        RECT  6.795 1.325 6.905 1.975 ;
        RECT  6.660 0.630 6.890 1.035 ;
        RECT  6.565 1.325 6.795 3.245 ;
        RECT  4.230 0.630 6.660 0.860 ;
        RECT  6.360 2.060 6.565 2.400 ;
        RECT  5.440 1.090 5.670 4.225 ;
        RECT  4.690 1.090 5.440 1.320 ;
        RECT  4.920 1.550 5.150 4.335 ;
        RECT  2.045 4.105 4.920 4.335 ;
        RECT  4.460 1.090 4.690 3.795 ;
        RECT  2.805 3.565 4.460 3.795 ;
        RECT  4.000 0.630 4.230 3.300 ;
        RECT  3.225 0.930 3.565 3.300 ;
        RECT  1.245 0.930 3.225 1.160 ;
        RECT  2.465 1.390 2.805 3.795 ;
        RECT  2.460 2.990 2.465 3.795 ;
        RECT  1.815 1.390 2.045 4.335 ;
        RECT  1.705 1.390 1.815 1.730 ;
        RECT  1.705 3.405 1.815 4.335 ;
        RECT  1.245 2.015 1.580 2.405 ;
        RECT  1.015 0.930 1.245 3.170 ;
        RECT  0.525 1.475 1.015 1.705 ;
        RECT  0.605 2.940 1.015 3.170 ;
        RECT  0.265 2.940 0.605 4.220 ;
        RECT  0.185 0.765 0.525 1.705 ;
    END
END AFHCINX2

MACRO CMPR42X2
    CLASS CORE ;
    FOREIGN CMPR42X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.400 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.185 0.765 26.220 1.575 ;
        RECT  26.185 2.380 26.220 3.555 ;
        RECT  25.955 0.765 26.185 3.555 ;
        RECT  25.880 0.765 25.955 1.575 ;
        RECT  25.880 2.380 25.955 3.555 ;
        END
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 0.945 0.520 1.755 ;
        RECT  0.400 2.745 0.520 3.555 ;
        RECT  0.180 0.945 0.400 3.555 ;
        RECT  0.170 1.235 0.180 3.265 ;
        END
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.895 1.875 23.045 2.105 ;
        RECT  22.665 1.285 22.895 2.105 ;
        RECT  22.655 1.285 22.665 1.515 ;
        END
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.945 1.985 17.470 2.215 ;
        RECT  16.715 1.845 16.945 2.240 ;
        RECT  15.060 2.010 16.715 2.240 ;
        RECT  14.830 2.010 15.060 2.665 ;
        RECT  14.620 2.435 14.830 2.665 ;
        END
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.730 2.965 20.905 3.195 ;
        RECT  20.520 1.265 20.730 3.360 ;
        RECT  20.500 1.265 20.520 3.445 ;
        RECT  20.115 1.265 20.500 1.495 ;
        RECT  20.180 3.105 20.500 3.445 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.195 4.175 17.250 4.405 ;
        RECT  16.285 4.175 17.195 4.410 ;
        RECT  16.055 4.085 16.285 4.410 ;
        RECT  14.405 4.085 16.055 4.315 ;
        RECT  14.175 4.005 14.405 4.315 ;
        RECT  13.375 4.005 14.175 4.235 ;
        RECT  13.145 4.005 13.375 4.410 ;
        RECT  10.425 4.180 13.145 4.410 ;
        RECT  10.195 4.005 10.425 4.410 ;
        RECT  9.390 4.005 10.195 4.235 ;
        RECT  9.160 4.005 9.390 4.405 ;
        RECT  7.060 4.175 9.160 4.405 ;
        RECT  6.830 4.005 7.060 4.405 ;
        RECT  4.175 4.005 6.830 4.235 ;
        RECT  3.895 4.005 4.175 4.340 ;
        RECT  3.665 4.005 3.895 4.410 ;
        RECT  3.350 4.180 3.665 4.410 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.010 2.525 8.450 2.755 ;
        RECT  7.780 2.525 8.010 2.985 ;
        RECT  6.565 2.755 7.780 2.985 ;
        RECT  6.335 2.755 6.565 3.625 ;
        RECT  5.295 3.395 6.335 3.625 ;
        RECT  5.295 2.265 5.350 2.495 ;
        RECT  5.065 2.265 5.295 3.625 ;
        RECT  3.820 2.265 5.065 2.495 ;
        RECT  3.440 2.265 3.820 2.635 ;
        RECT  2.070 2.265 3.440 2.495 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.800 6.515 2.030 ;
        RECT  1.690 1.800 1.765 2.075 ;
        RECT  1.535 1.800 1.690 2.415 ;
        RECT  1.460 1.845 1.535 2.415 ;
        RECT  1.245 2.185 1.460 2.415 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.460 -0.400 26.400 0.400 ;
        RECT  25.120 -0.400 25.460 0.575 ;
        RECT  22.655 -0.400 25.120 0.400 ;
        RECT  22.315 -0.400 22.655 0.575 ;
        RECT  21.450 -0.400 22.315 0.400 ;
        RECT  21.110 -0.400 21.450 0.575 ;
        RECT  17.315 -0.400 21.110 0.400 ;
        RECT  16.975 -0.400 17.315 0.575 ;
        RECT  13.205 -0.400 16.975 0.400 ;
        RECT  12.865 -0.400 13.205 0.575 ;
        RECT  9.650 -0.400 12.865 0.400 ;
        RECT  9.310 -0.400 9.650 0.575 ;
        RECT  6.850 -0.400 9.310 0.400 ;
        RECT  6.510 -0.400 6.850 0.575 ;
        RECT  5.380 -0.400 6.510 0.400 ;
        RECT  5.040 -0.400 5.380 0.575 ;
        RECT  3.860 -0.400 5.040 0.400 ;
        RECT  3.520 -0.400 3.860 0.575 ;
        RECT  1.280 -0.400 3.520 0.400 ;
        RECT  0.940 -0.400 1.280 0.575 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  25.460 4.640 26.400 5.440 ;
        RECT  25.405 4.465 25.460 5.440 ;
        RECT  25.175 3.320 25.405 5.440 ;
        RECT  25.120 4.465 25.175 5.440 ;
        RECT  22.405 4.640 25.120 5.440 ;
        RECT  22.065 4.465 22.405 5.440 ;
        RECT  17.710 4.640 22.065 5.440 ;
        RECT  17.480 3.710 17.710 5.440 ;
        RECT  17.250 3.710 17.480 3.940 ;
        RECT  13.945 4.640 17.480 5.440 ;
        RECT  16.910 3.130 17.250 3.940 ;
        RECT  13.605 4.465 13.945 5.440 ;
        RECT  9.960 4.640 13.605 5.440 ;
        RECT  9.620 4.465 9.960 5.440 ;
        RECT  6.600 4.640 9.620 5.440 ;
        RECT  6.260 4.465 6.600 5.440 ;
        RECT  5.540 4.640 6.260 5.440 ;
        RECT  5.200 4.465 5.540 5.440 ;
        RECT  1.280 4.640 5.200 5.440 ;
        RECT  0.940 3.840 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  25.430 1.920 25.725 2.150 ;
        RECT  25.200 0.805 25.430 3.090 ;
        RECT  23.795 0.805 25.200 1.035 ;
        RECT  24.945 2.860 25.200 3.090 ;
        RECT  24.740 1.265 24.970 2.630 ;
        RECT  24.890 2.860 24.945 4.190 ;
        RECT  24.715 2.860 24.890 4.250 ;
        RECT  23.550 1.265 24.740 1.495 ;
        RECT  24.485 2.400 24.740 2.630 ;
        RECT  24.660 3.960 24.715 4.250 ;
        RECT  23.885 4.020 24.660 4.250 ;
        RECT  23.505 1.725 24.510 1.955 ;
        RECT  24.430 2.400 24.485 3.405 ;
        RECT  24.255 2.400 24.430 3.790 ;
        RECT  24.200 3.175 24.255 3.790 ;
        RECT  23.165 3.560 24.200 3.790 ;
        RECT  23.970 2.580 24.025 2.945 ;
        RECT  23.795 2.580 23.970 3.330 ;
        RECT  23.545 4.020 23.885 4.360 ;
        RECT  23.740 2.715 23.795 3.330 ;
        RECT  21.835 3.100 23.740 3.330 ;
        RECT  23.320 0.800 23.550 1.495 ;
        RECT  23.275 1.725 23.505 2.775 ;
        RECT  23.075 0.800 23.320 1.030 ;
        RECT  22.350 2.545 23.275 2.775 ;
        RECT  23.055 3.560 23.165 3.920 ;
        RECT  22.880 3.560 23.055 4.235 ;
        RECT  22.825 3.580 22.880 4.235 ;
        RECT  21.650 4.005 22.825 4.235 ;
        RECT  22.120 0.805 22.350 2.775 ;
        RECT  21.250 0.805 22.120 1.035 ;
        RECT  21.820 1.430 21.835 3.330 ;
        RECT  21.730 1.375 21.820 3.330 ;
        RECT  21.605 1.375 21.730 3.685 ;
        RECT  21.420 4.005 21.650 4.410 ;
        RECT  21.480 1.375 21.605 1.715 ;
        RECT  21.500 2.795 21.605 3.685 ;
        RECT  21.190 3.455 21.500 3.685 ;
        RECT  19.580 4.180 21.420 4.410 ;
        RECT  21.250 1.945 21.375 2.370 ;
        RECT  21.145 0.805 21.250 2.370 ;
        RECT  20.960 3.455 21.190 3.950 ;
        RECT  21.020 0.805 21.145 2.175 ;
        RECT  20.370 0.805 21.020 1.035 ;
        RECT  19.810 3.720 20.960 3.950 ;
        RECT  20.140 0.630 20.370 1.035 ;
        RECT  20.040 1.725 20.270 2.875 ;
        RECT  18.480 0.630 20.140 0.860 ;
        RECT  19.715 1.725 20.040 1.955 ;
        RECT  19.780 2.645 20.040 2.875 ;
        RECT  19.115 2.185 19.810 2.415 ;
        RECT  19.580 2.645 19.780 3.475 ;
        RECT  19.485 1.130 19.715 1.955 ;
        RECT  19.550 2.645 19.580 4.410 ;
        RECT  19.440 3.135 19.550 4.410 ;
        RECT  19.375 1.130 19.485 1.470 ;
        RECT  19.350 3.245 19.440 4.410 ;
        RECT  19.060 2.000 19.115 3.395 ;
        RECT  18.940 2.000 19.060 3.975 ;
        RECT  18.885 1.105 18.940 3.975 ;
        RECT  18.710 1.105 18.885 2.230 ;
        RECT  18.720 3.165 18.885 3.975 ;
        RECT  18.480 2.505 18.655 2.920 ;
        RECT  18.425 0.630 18.480 2.920 ;
        RECT  18.250 0.630 18.425 2.735 ;
        RECT  18.000 3.160 18.340 3.970 ;
        RECT  18.180 0.630 18.250 1.035 ;
        RECT  16.580 0.805 18.180 1.035 ;
        RECT  17.950 1.265 18.020 1.985 ;
        RECT  17.950 3.160 18.000 3.390 ;
        RECT  17.790 1.265 17.950 3.390 ;
        RECT  17.720 1.755 17.790 3.390 ;
        RECT  17.650 2.470 17.720 3.390 ;
        RECT  15.290 2.470 17.650 2.700 ;
        RECT  16.350 0.630 16.580 1.035 ;
        RECT  16.290 1.270 16.555 1.500 ;
        RECT  13.680 0.630 16.350 0.860 ;
        RECT  16.060 1.270 16.290 1.780 ;
        RECT  14.225 3.085 16.160 3.315 ;
        RECT  14.600 1.550 16.060 1.780 ;
        RECT  14.140 1.090 15.735 1.320 ;
        RECT  13.700 3.545 15.440 3.775 ;
        RECT  14.370 1.550 14.600 1.955 ;
        RECT  14.325 1.725 14.370 1.955 ;
        RECT  14.225 1.725 14.325 2.400 ;
        RECT  14.095 1.725 14.225 3.315 ;
        RECT  13.910 1.090 14.140 1.495 ;
        RECT  13.995 2.115 14.095 3.315 ;
        RECT  13.885 2.115 13.995 2.455 ;
        RECT  12.455 1.265 13.910 1.495 ;
        RECT  13.470 3.005 13.700 3.775 ;
        RECT  13.450 0.630 13.680 1.035 ;
        RECT  12.710 3.005 13.470 3.235 ;
        RECT  11.985 0.805 13.450 1.035 ;
        RECT  12.915 3.465 13.240 3.695 ;
        RECT  12.685 3.465 12.915 3.950 ;
        RECT  12.455 2.890 12.710 3.235 ;
        RECT  10.885 3.720 12.685 3.950 ;
        RECT  12.225 1.265 12.455 3.490 ;
        RECT  12.215 1.265 12.225 1.625 ;
        RECT  11.350 3.260 12.225 3.490 ;
        RECT  11.985 1.980 11.995 3.030 ;
        RECT  11.765 0.805 11.985 3.030 ;
        RECT  11.755 0.805 11.765 2.210 ;
        RECT  11.645 2.800 11.765 3.030 ;
        RECT  11.315 1.210 11.755 1.495 ;
        RECT  11.295 1.745 11.525 2.120 ;
        RECT  11.120 2.560 11.350 3.490 ;
        RECT  10.975 1.155 11.315 1.495 ;
        RECT  10.460 1.745 11.295 1.975 ;
        RECT  10.855 2.560 11.120 2.790 ;
        RECT  10.655 3.545 10.885 3.950 ;
        RECT  10.625 2.210 10.855 2.790 ;
        RECT  10.340 3.020 10.725 3.250 ;
        RECT  9.745 3.545 10.655 3.775 ;
        RECT  10.340 1.155 10.460 1.975 ;
        RECT  10.120 1.155 10.340 3.250 ;
        RECT  10.110 1.210 10.120 3.250 ;
        RECT  9.515 0.935 9.745 3.775 ;
        RECT  8.330 0.935 9.515 1.165 ;
        RECT  8.930 3.545 9.515 3.775 ;
        RECT  8.930 1.395 9.160 2.765 ;
        RECT  7.610 1.395 8.930 1.625 ;
        RECT  8.910 2.535 8.930 2.765 ;
        RECT  8.700 3.545 8.930 3.945 ;
        RECT  8.680 2.535 8.910 3.240 ;
        RECT  7.550 1.855 8.700 2.085 ;
        RECT  7.740 3.715 8.700 3.945 ;
        RECT  8.470 3.010 8.680 3.240 ;
        RECT  8.240 3.010 8.470 3.485 ;
        RECT  7.990 0.825 8.330 1.165 ;
        RECT  7.020 3.255 8.240 3.485 ;
        RECT  7.380 1.020 7.610 1.625 ;
        RECT  7.320 1.855 7.550 2.525 ;
        RECT  7.270 1.020 7.380 1.360 ;
        RECT  6.975 2.295 7.320 2.525 ;
        RECT  6.745 1.340 6.975 2.525 ;
        RECT  5.980 1.340 6.745 1.570 ;
        RECT  6.100 2.295 6.745 2.525 ;
        RECT  5.870 2.295 6.100 3.155 ;
        RECT  5.745 1.120 5.980 1.570 ;
        RECT  5.760 2.815 5.870 3.155 ;
        RECT  5.640 1.120 5.745 1.460 ;
        RECT  4.440 2.875 4.780 3.685 ;
        RECT  4.565 0.865 4.620 1.205 ;
        RECT  4.280 0.865 4.565 1.320 ;
        RECT  3.320 3.380 4.440 3.610 ;
        RECT  3.320 1.090 4.280 1.320 ;
        RECT  3.035 1.090 3.320 1.570 ;
        RECT  2.980 3.325 3.320 3.665 ;
        RECT  2.980 1.230 3.035 1.570 ;
        RECT  2.260 1.150 2.600 1.490 ;
        RECT  2.260 3.325 2.600 3.665 ;
        RECT  0.980 1.205 2.260 1.435 ;
        RECT  0.980 3.380 2.260 3.610 ;
        RECT  0.750 1.205 0.980 3.610 ;
        RECT  0.630 2.175 0.750 2.515 ;
    END
END CMPR42X2

MACRO CMPR42X1
    CLASS CORE ;
    FOREIGN CMPR42X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CMPR42X2 ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.220 1.175 22.265 3.265 ;
        RECT  22.035 1.120 22.220 3.555 ;
        RECT  21.880 1.120 22.035 1.460 ;
        RECT  21.920 2.380 22.035 3.555 ;
        RECT  21.880 2.745 21.920 3.555 ;
        END
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 1.355 0.520 1.695 ;
        RECT  0.400 2.745 0.520 3.555 ;
        RECT  0.180 1.355 0.400 3.555 ;
        RECT  0.170 1.410 0.180 3.265 ;
        END
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.055 2.375 19.585 2.660 ;
        RECT  18.715 2.320 19.055 2.660 ;
        END
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.340 1.800 14.000 2.140 ;
        RECT  12.845 1.800 13.340 2.030 ;
        RECT  12.615 1.590 12.845 2.030 ;
        END
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.940 1.370 16.995 1.845 ;
        RECT  16.945 2.635 16.995 3.080 ;
        RECT  16.940 2.635 16.945 3.195 ;
        RECT  16.715 1.370 16.940 3.195 ;
        RECT  16.710 1.370 16.715 3.080 ;
        RECT  16.655 1.370 16.710 1.845 ;
        RECT  16.655 2.635 16.710 3.080 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.060 3.950 13.090 4.290 ;
        RECT  12.750 3.500 13.060 4.290 ;
        RECT  12.680 3.500 12.750 4.235 ;
        RECT  6.305 4.005 12.680 4.235 ;
        RECT  6.075 4.005 6.305 4.410 ;
        RECT  3.030 4.180 6.075 4.410 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.880 3.990 2.110 ;
        RECT  3.515 1.845 3.745 2.110 ;
        RECT  2.100 1.880 3.515 2.110 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.650 1.985 4.760 2.325 ;
        RECT  4.420 1.985 4.650 2.570 ;
        RECT  1.765 2.340 4.420 2.570 ;
        RECT  1.535 1.845 1.765 2.570 ;
        RECT  1.300 2.100 1.535 2.440 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.420 -0.400 22.440 0.400 ;
        RECT  21.080 -0.400 21.420 0.575 ;
        RECT  18.225 -0.400 21.080 0.400 ;
        RECT  17.415 -0.400 18.225 0.575 ;
        RECT  13.850 -0.400 17.415 0.400 ;
        RECT  13.510 -0.400 13.850 0.575 ;
        RECT  10.660 -0.400 13.510 0.400 ;
        RECT  10.320 -0.400 10.660 0.575 ;
        RECT  7.780 -0.400 10.320 0.400 ;
        RECT  7.440 -0.400 7.780 0.575 ;
        RECT  5.020 -0.400 7.440 0.400 ;
        RECT  4.680 -0.400 5.020 1.275 ;
        RECT  2.720 -0.400 4.680 0.400 ;
        RECT  2.380 -0.400 2.720 0.575 ;
        RECT  1.120 -0.400 2.380 0.400 ;
        RECT  0.780 -0.400 1.120 0.575 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.655 4.640 22.440 5.440 ;
        RECT  21.315 4.465 21.655 5.440 ;
        RECT  18.775 4.640 21.315 5.440 ;
        RECT  18.435 3.810 18.775 5.440 ;
        RECT  17.755 4.640 18.435 5.440 ;
        RECT  17.415 4.465 17.755 5.440 ;
        RECT  13.660 4.640 17.415 5.440 ;
        RECT  13.320 2.885 13.660 5.440 ;
        RECT  11.060 4.640 13.320 5.440 ;
        RECT  10.720 4.465 11.060 5.440 ;
        RECT  7.580 4.640 10.720 5.440 ;
        RECT  7.240 4.465 7.580 5.440 ;
        RECT  2.800 4.640 7.240 5.440 ;
        RECT  4.925 3.410 4.980 3.750 ;
        RECT  4.640 3.410 4.925 3.950 ;
        RECT  2.800 3.720 4.640 3.950 ;
        RECT  2.570 3.720 2.800 5.440 ;
        RECT  2.460 4.465 2.570 5.440 ;
        RECT  1.280 4.640 2.460 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.650 1.805 21.805 2.145 ;
        RECT  21.420 1.555 21.650 4.040 ;
        RECT  20.795 1.555 21.420 1.785 ;
        RECT  20.295 3.810 21.420 4.040 ;
        RECT  20.980 2.015 21.135 2.355 ;
        RECT  20.750 2.015 20.980 3.580 ;
        RECT  20.565 0.785 20.795 1.785 ;
        RECT  20.320 2.015 20.750 2.245 ;
        RECT  19.535 3.350 20.750 3.580 ;
        RECT  19.720 0.785 20.565 1.015 ;
        RECT  20.180 2.780 20.520 3.120 ;
        RECT  20.090 1.245 20.320 2.245 ;
        RECT  19.955 3.810 20.295 4.150 ;
        RECT  18.365 2.890 20.180 3.120 ;
        RECT  19.260 1.245 20.090 1.475 ;
        RECT  18.365 1.705 19.610 1.935 ;
        RECT  19.195 3.350 19.535 3.790 ;
        RECT  19.030 0.760 19.260 1.475 ;
        RECT  17.955 3.350 19.195 3.580 ;
        RECT  18.920 0.760 19.030 1.100 ;
        RECT  18.135 1.375 18.365 3.120 ;
        RECT  18.015 1.375 18.135 1.715 ;
        RECT  18.015 2.740 18.135 3.120 ;
        RECT  17.480 2.890 18.015 3.120 ;
        RECT  17.725 3.350 17.955 4.145 ;
        RECT  17.785 2.030 17.905 2.370 ;
        RECT  17.555 0.805 17.785 2.370 ;
        RECT  17.075 3.915 17.725 4.145 ;
        RECT  17.050 0.805 17.555 1.035 ;
        RECT  17.250 2.890 17.480 3.685 ;
        RECT  16.615 3.455 17.250 3.685 ;
        RECT  16.845 3.915 17.075 4.380 ;
        RECT  16.820 0.630 17.050 1.035 ;
        RECT  15.895 4.150 16.845 4.380 ;
        RECT  14.920 0.630 16.820 0.860 ;
        RECT  16.385 3.455 16.615 3.920 ;
        RECT  16.125 3.690 16.385 3.920 ;
        RECT  16.035 1.105 16.235 1.445 ;
        RECT  15.895 1.105 16.035 3.225 ;
        RECT  15.805 1.105 15.895 4.380 ;
        RECT  15.665 2.885 15.805 4.380 ;
        RECT  15.380 4.065 15.435 4.405 ;
        RECT  15.150 1.105 15.380 4.405 ;
        RECT  14.975 2.955 15.150 3.295 ;
        RECT  15.095 4.065 15.150 4.405 ;
        RECT  14.690 0.630 14.920 2.695 ;
        RECT  13.280 0.805 14.690 1.035 ;
        RECT  14.420 1.320 14.460 2.600 ;
        RECT  14.230 1.320 14.420 3.295 ;
        RECT  14.120 1.320 14.230 1.550 ;
        RECT  14.080 2.370 14.230 3.295 ;
        RECT  12.660 2.370 14.080 2.600 ;
        RECT  13.050 0.630 13.280 1.035 ;
        RECT  11.145 0.630 13.050 0.860 ;
        RECT  12.560 2.830 12.900 3.170 ;
        RECT  12.385 1.090 12.820 1.320 ;
        RECT  12.320 2.260 12.660 2.600 ;
        RECT  11.180 2.830 12.560 3.060 ;
        RECT  12.155 1.090 12.385 1.955 ;
        RECT  11.840 3.295 12.180 3.635 ;
        RECT  11.180 1.725 12.155 1.955 ;
        RECT  11.695 1.090 11.925 1.495 ;
        RECT  10.360 3.295 11.840 3.525 ;
        RECT  10.385 1.265 11.695 1.495 ;
        RECT  10.950 1.725 11.180 3.060 ;
        RECT  10.915 0.630 11.145 1.035 ;
        RECT  10.840 2.260 10.950 2.600 ;
        RECT  9.530 0.805 10.915 1.035 ;
        RECT  10.385 1.890 10.440 2.230 ;
        RECT  10.360 1.265 10.385 2.230 ;
        RECT  10.155 1.265 10.360 3.695 ;
        RECT  9.820 1.265 10.155 1.495 ;
        RECT  10.130 1.890 10.155 3.695 ;
        RECT  10.100 1.890 10.130 2.230 ;
        RECT  10.020 2.885 10.130 3.695 ;
        RECT  9.530 2.885 9.640 3.695 ;
        RECT  9.300 0.805 9.530 3.695 ;
        RECT  9.100 1.155 9.300 1.495 ;
        RECT  7.775 3.545 8.880 3.775 ;
        RECT  8.530 1.155 8.575 1.495 ;
        RECT  8.390 0.630 8.530 1.495 ;
        RECT  8.345 0.630 8.390 3.075 ;
        RECT  8.190 0.630 8.345 3.130 ;
        RECT  8.160 1.210 8.190 3.130 ;
        RECT  8.005 2.790 8.160 3.130 ;
        RECT  7.775 2.220 7.930 2.560 ;
        RECT  7.545 1.090 7.775 3.775 ;
        RECT  6.460 1.090 7.545 1.320 ;
        RECT  6.460 3.545 7.545 3.775 ;
        RECT  7.150 1.985 7.260 2.325 ;
        RECT  6.920 1.775 7.150 3.060 ;
        RECT  5.740 1.775 6.920 2.005 ;
        RECT  5.685 2.830 6.920 3.060 ;
        RECT  6.120 0.980 6.460 1.320 ;
        RECT  6.175 3.295 6.460 3.775 ;
        RECT  6.120 3.295 6.175 3.635 ;
        RECT  5.640 2.260 5.980 2.600 ;
        RECT  5.510 0.955 5.740 2.005 ;
        RECT  5.455 2.830 5.685 3.675 ;
        RECT  5.220 2.315 5.640 2.600 ;
        RECT  5.400 0.955 5.510 1.295 ;
        RECT  4.990 1.525 5.220 3.160 ;
        RECT  4.450 1.525 4.990 1.755 ;
        RECT  4.180 2.930 4.990 3.160 ;
        RECT  4.220 1.145 4.450 1.755 ;
        RECT  3.880 1.035 4.220 1.375 ;
        RECT  3.840 2.930 4.180 3.275 ;
        RECT  3.410 1.235 3.520 1.575 ;
        RECT  3.370 2.920 3.480 3.260 ;
        RECT  3.180 0.805 3.410 1.575 ;
        RECT  3.140 2.920 3.370 3.490 ;
        RECT  1.920 0.805 3.180 1.035 ;
        RECT  2.040 3.260 3.140 3.490 ;
        RECT  0.980 2.800 2.760 3.030 ;
        RECT  2.380 1.295 2.720 1.635 ;
        RECT  0.980 1.350 2.380 1.580 ;
        RECT  1.810 3.260 2.040 4.345 ;
        RECT  1.635 0.630 1.920 1.035 ;
        RECT  1.700 4.005 1.810 4.345 ;
        RECT  1.580 0.630 1.635 0.970 ;
        RECT  0.750 1.350 0.980 3.030 ;
        RECT  0.630 2.030 0.750 2.370 ;
    END
END CMPR42X1

MACRO CMPR32X1
    CLASS CORE ;
    FOREIGN CMPR32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.570 1.285 13.645 1.515 ;
        RECT  13.460 1.285 13.570 1.845 ;
        RECT  13.460 2.635 13.570 3.605 ;
        RECT  13.230 1.285 13.460 3.605 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.005 2.380 12.325 2.660 ;
        RECT  11.985 1.430 12.005 2.660 ;
        RECT  11.755 1.430 11.985 3.135 ;
        RECT  11.665 1.430 11.755 1.770 ;
        RECT  11.645 2.795 11.755 3.135 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.220 1.820 9.485 2.050 ;
        RECT  8.990 1.820 9.220 3.220 ;
        RECT  8.600 2.865 8.990 3.220 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.040 0.760 2.380 ;
        RECT  0.420 2.040 0.445 2.635 ;
        RECT  0.215 2.150 0.420 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.895 2.350 4.835 2.690 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.770 -0.400 13.860 0.400 ;
        RECT  12.430 -0.400 12.770 1.615 ;
        RECT  10.080 -0.400 12.430 0.400 ;
        RECT  9.740 -0.400 10.080 0.575 ;
        RECT  4.725 -0.400 9.740 0.400 ;
        RECT  4.385 -0.400 4.725 0.900 ;
        RECT  1.285 -0.400 4.385 0.400 ;
        RECT  0.945 -0.400 1.285 0.575 ;
        RECT  0.000 -0.400 0.945 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.775 4.640 13.860 5.440 ;
        RECT  12.435 3.930 12.775 5.440 ;
        RECT  8.935 4.640 12.435 5.440 ;
        RECT  8.595 4.465 8.935 5.440 ;
        RECT  1.200 4.640 8.595 5.440 ;
        RECT  0.860 4.465 1.200 5.440 ;
        RECT  0.000 4.640 0.860 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.635 2.015 12.865 3.595 ;
        RECT  11.645 3.365 12.635 3.595 ;
        RECT  11.415 3.365 11.645 3.945 ;
        RECT  9.395 4.180 11.455 4.410 ;
        RECT  10.455 3.715 11.415 3.945 ;
        RECT  11.140 0.630 11.295 0.860 ;
        RECT  11.140 3.120 11.175 3.460 ;
        RECT  10.910 0.630 11.140 3.460 ;
        RECT  10.900 0.630 10.910 1.040 ;
        RECT  10.835 3.120 10.910 3.460 ;
        RECT  9.495 0.810 10.900 1.040 ;
        RECT  10.455 1.345 10.680 1.770 ;
        RECT  10.450 1.345 10.455 3.945 ;
        RECT  10.225 1.540 10.450 3.945 ;
        RECT  10.115 3.215 10.225 3.555 ;
        RECT  9.730 1.270 9.960 2.875 ;
        RECT  9.035 1.270 9.730 1.500 ;
        RECT  9.680 2.645 9.730 2.875 ;
        RECT  9.450 2.645 9.680 3.555 ;
        RECT  9.265 0.630 9.495 1.040 ;
        RECT  9.165 4.005 9.395 4.410 ;
        RECT  5.880 0.630 9.265 0.860 ;
        RECT  7.855 4.005 9.165 4.235 ;
        RECT  8.805 1.090 9.035 1.500 ;
        RECT  6.670 1.090 8.805 1.320 ;
        RECT  8.570 2.195 8.760 2.535 ;
        RECT  8.340 1.585 8.570 2.535 ;
        RECT  8.315 2.305 8.340 2.535 ;
        RECT  8.085 2.305 8.315 3.770 ;
        RECT  7.850 3.580 7.855 4.235 ;
        RECT  7.625 1.585 7.850 4.235 ;
        RECT  7.620 1.585 7.625 3.810 ;
        RECT  7.175 3.580 7.620 3.810 ;
        RECT  7.160 1.790 7.390 3.350 ;
        RECT  7.130 1.790 7.160 2.020 ;
        RECT  6.795 3.120 7.160 3.350 ;
        RECT  6.900 1.585 7.130 2.020 ;
        RECT  6.670 2.360 6.930 2.700 ;
        RECT  6.685 3.120 6.795 3.780 ;
        RECT  6.565 3.120 6.685 4.410 ;
        RECT  6.440 1.090 6.670 2.890 ;
        RECT  6.455 3.440 6.565 4.410 ;
        RECT  5.255 4.055 6.455 4.410 ;
        RECT  6.175 2.655 6.440 2.890 ;
        RECT  5.300 2.070 6.210 2.420 ;
        RECT  6.075 2.655 6.175 3.425 ;
        RECT  5.945 2.655 6.075 3.480 ;
        RECT  5.765 3.140 5.945 3.480 ;
        RECT  5.650 0.630 5.880 1.750 ;
        RECT  5.735 3.140 5.765 3.825 ;
        RECT  5.535 3.195 5.735 3.825 ;
        RECT  5.540 1.135 5.650 1.750 ;
        RECT  4.155 1.135 5.540 1.365 ;
        RECT  3.440 3.595 5.535 3.825 ;
        RECT  5.070 1.635 5.300 3.365 ;
        RECT  1.660 4.180 5.255 4.410 ;
        RECT  3.695 1.635 5.070 1.865 ;
        RECT  3.900 3.135 5.070 3.365 ;
        RECT  3.925 0.875 4.155 1.365 ;
        RECT  2.450 0.875 3.925 1.105 ;
        RECT  3.670 2.980 3.900 3.365 ;
        RECT  3.465 1.440 3.695 1.865 ;
        RECT  3.210 3.030 3.440 3.825 ;
        RECT  3.180 3.030 3.210 3.260 ;
        RECT  2.950 2.075 3.180 3.260 ;
        RECT  2.750 3.495 2.980 3.950 ;
        RECT  2.910 2.075 2.950 2.305 ;
        RECT  2.680 1.420 2.910 2.305 ;
        RECT  2.125 3.495 2.750 3.725 ;
        RECT  2.450 2.535 2.620 3.265 ;
        RECT  2.390 0.875 2.450 3.265 ;
        RECT  2.220 0.875 2.390 2.765 ;
        RECT  1.990 3.050 2.125 3.725 ;
        RECT  1.895 1.395 1.990 3.725 ;
        RECT  1.760 1.395 1.895 3.280 ;
        RECT  1.505 2.940 1.760 3.280 ;
        RECT  1.430 3.655 1.660 4.410 ;
        RECT  1.380 2.040 1.490 2.380 ;
        RECT  1.235 3.655 1.430 3.885 ;
        RECT  1.235 1.395 1.380 2.380 ;
        RECT  1.150 1.395 1.235 3.885 ;
        RECT  0.520 1.395 1.150 1.625 ;
        RECT  1.005 2.095 1.150 3.885 ;
        RECT  0.180 2.890 1.005 3.230 ;
        RECT  0.180 0.815 0.520 1.625 ;
    END
END CMPR32X1

MACRO CMPR22X1
    CLASS CORE ;
    FOREIGN CMPR22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.330 4.235 3.220 ;
        RECT  3.590 1.330 4.005 1.560 ;
        RECT  3.245 2.840 4.005 3.220 ;
        RECT  3.360 1.210 3.590 1.560 ;
        RECT  3.015 2.840 3.245 3.730 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.610 1.845 7.705 2.075 ;
        RECT  7.400 1.380 7.610 2.075 ;
        RECT  7.380 1.380 7.400 3.115 ;
        RECT  7.185 1.845 7.380 3.115 ;
        RECT  7.170 1.845 7.185 3.970 ;
        RECT  6.955 2.885 7.170 3.970 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 2.520 6.065 3.445 ;
        RECT  5.160 3.215 5.835 3.445 ;
        RECT  4.930 3.215 5.160 4.235 ;
        RECT  2.785 4.005 4.930 4.235 ;
        RECT  3.545 1.800 3.775 2.520 ;
        RECT  2.785 2.290 3.545 2.520 ;
        RECT  2.555 2.290 2.785 4.235 ;
        RECT  2.195 2.290 2.555 2.660 ;
        RECT  2.115 2.290 2.195 2.575 ;
        RECT  1.775 2.235 2.115 2.575 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.820 5.075 2.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.150 -0.400 7.920 0.400 ;
        RECT  6.920 -0.400 7.150 1.355 ;
        RECT  5.125 -0.400 6.920 0.400 ;
        RECT  6.815 1.125 6.920 1.355 ;
        RECT  6.585 1.125 6.815 1.720 ;
        RECT  4.785 -0.400 5.125 0.575 ;
        RECT  1.360 -0.400 4.785 0.400 ;
        RECT  1.020 -0.400 1.360 0.575 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.480 4.640 7.920 5.440 ;
        RECT  6.140 4.465 6.480 5.440 ;
        RECT  4.780 4.640 6.140 5.440 ;
        RECT  4.440 4.465 4.780 5.440 ;
        RECT  1.280 4.640 4.440 5.440 ;
        RECT  0.940 4.465 1.280 5.440 ;
        RECT  0.000 4.640 0.940 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.525 1.980 6.840 2.320 ;
        RECT  6.350 0.665 6.690 0.895 ;
        RECT  6.350 1.980 6.525 3.905 ;
        RECT  6.295 0.665 6.350 3.905 ;
        RECT  6.120 0.665 6.295 2.210 ;
        RECT  5.625 3.675 6.295 3.905 ;
        RECT  5.600 1.210 5.885 1.550 ;
        RECT  5.395 3.675 5.625 4.085 ;
        RECT  5.545 1.210 5.600 2.985 ;
        RECT  5.370 1.265 5.545 2.985 ;
        RECT  4.700 1.265 5.370 1.495 ;
        RECT  4.700 2.755 5.370 2.985 ;
        RECT  4.470 0.805 4.700 1.495 ;
        RECT  4.470 2.755 4.700 3.775 ;
        RECT  4.365 0.805 4.470 1.035 ;
        RECT  3.680 3.545 4.470 3.775 ;
        RECT  4.025 0.675 4.365 1.035 ;
        RECT  3.130 0.675 4.025 0.905 ;
        RECT  2.900 0.675 3.130 1.955 ;
        RECT  1.385 1.725 2.900 1.955 ;
        RECT  2.440 0.630 2.670 1.035 ;
        RECT  0.925 1.265 2.550 1.495 ;
        RECT  0.465 0.805 2.440 1.035 ;
        RECT  2.095 4.005 2.325 4.405 ;
        RECT  0.465 4.005 2.095 4.235 ;
        RECT  1.500 3.180 1.840 3.520 ;
        RECT  0.925 3.180 1.500 3.410 ;
        RECT  1.155 1.725 1.385 2.560 ;
        RECT  0.695 1.265 0.925 3.410 ;
        RECT  0.235 0.760 0.465 4.235 ;
    END
END CMPR22X1

MACRO BMXX1
    CLASS CORE ;
    FOREIGN BMXX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 2.160 9.840 2.715 ;
        END
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.690 2.185 7.120 2.665 ;
        END
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.305 2.635 12.360 3.635 ;
        RECT  12.075 1.265 12.305 3.635 ;
        RECT  12.020 2.825 12.075 3.635 ;
        END
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.930 1.790 6.460 2.270 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.820 1.110 2.540 ;
        RECT  0.770 2.200 0.800 2.540 ;
        END
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 2.010 1.800 2.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.360 -0.400 12.540 0.400 ;
        RECT  12.020 -0.400 12.360 0.575 ;
        RECT  8.625 -0.400 12.020 0.400 ;
        RECT  8.285 -0.400 8.625 0.575 ;
        RECT  6.605 -0.400 8.285 0.400 ;
        RECT  6.265 -0.400 6.605 0.575 ;
        RECT  1.320 -0.400 6.265 0.400 ;
        RECT  0.980 -0.400 1.320 1.520 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.935 4.640 12.540 5.440 ;
        RECT  11.595 4.465 11.935 5.440 ;
        RECT  9.090 4.640 11.595 5.440 ;
        RECT  6.400 4.465 9.090 5.440 ;
        RECT  1.320 4.640 6.400 5.440 ;
        RECT  0.980 3.920 1.320 5.440 ;
        RECT  0.000 4.640 0.980 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.790 1.085 11.805 2.595 ;
        RECT  11.575 0.665 11.790 2.595 ;
        RECT  11.560 0.665 11.575 1.315 ;
        RECT  11.515 2.365 11.575 2.595 ;
        RECT  10.960 0.665 11.560 0.895 ;
        RECT  11.365 2.365 11.515 3.985 ;
        RECT  11.285 2.365 11.365 4.375 ;
        RECT  11.330 1.650 11.345 2.135 ;
        RECT  11.115 1.125 11.330 2.135 ;
        RECT  11.135 3.755 11.285 4.375 ;
        RECT  9.665 4.145 11.135 4.375 ;
        RECT  11.100 1.125 11.115 1.880 ;
        RECT  10.300 1.125 11.100 1.355 ;
        RECT  10.620 0.630 10.960 0.895 ;
        RECT  10.905 2.855 10.915 3.365 ;
        RECT  10.870 2.855 10.905 3.810 ;
        RECT  10.675 1.585 10.870 3.810 ;
        RECT  10.640 1.585 10.675 3.085 ;
        RECT  8.690 3.580 10.675 3.810 ;
        RECT  10.530 1.585 10.640 1.815 ;
        RECT  9.535 0.630 10.620 0.860 ;
        RECT  10.070 1.125 10.300 3.320 ;
        RECT  9.770 1.460 10.070 1.690 ;
        RECT  9.865 3.090 10.070 3.320 ;
        RECT  9.150 3.060 9.445 3.290 ;
        RECT  9.150 1.430 9.335 1.930 ;
        RECT  5.980 0.805 9.195 1.035 ;
        RECT  9.105 1.430 9.150 3.290 ;
        RECT  8.920 1.700 9.105 3.290 ;
        RECT  8.460 2.995 8.690 3.810 ;
        RECT  8.070 2.995 8.460 3.225 ;
        RECT  7.840 1.265 8.070 3.225 ;
        RECT  7.830 3.695 7.980 3.925 ;
        RECT  7.725 1.265 7.840 1.495 ;
        RECT  7.600 3.695 7.830 4.235 ;
        RECT  5.900 4.005 7.600 4.235 ;
        RECT  7.370 1.725 7.580 3.195 ;
        RECT  7.365 1.725 7.370 3.775 ;
        RECT  7.350 1.265 7.365 3.775 ;
        RECT  7.135 1.265 7.350 1.955 ;
        RECT  7.140 2.965 7.350 3.775 ;
        RECT  5.440 3.545 7.140 3.775 ;
        RECT  7.025 1.265 7.135 1.605 ;
        RECT  5.750 0.630 5.980 1.035 ;
        RECT  5.700 2.830 5.980 3.170 ;
        RECT  5.670 4.005 5.900 4.405 ;
        RECT  5.700 1.330 5.875 1.560 ;
        RECT  4.400 0.630 5.750 0.860 ;
        RECT  5.640 1.330 5.700 3.170 ;
        RECT  3.020 4.175 5.670 4.405 ;
        RECT  5.470 1.330 5.640 3.115 ;
        RECT  5.210 2.210 5.470 2.550 ;
        RECT  5.210 3.545 5.440 3.945 ;
        RECT  4.970 2.850 5.240 3.190 ;
        RECT  3.480 3.715 5.210 3.945 ;
        RECT  4.970 1.090 5.175 1.320 ;
        RECT  4.740 1.090 4.970 3.485 ;
        RECT  3.940 3.255 4.740 3.485 ;
        RECT  4.400 2.795 4.510 3.025 ;
        RECT  4.170 0.630 4.400 3.025 ;
        RECT  3.710 0.630 3.940 3.485 ;
        RECT  2.040 0.630 3.710 0.860 ;
        RECT  3.250 1.090 3.480 3.945 ;
        RECT  3.140 1.090 3.250 1.320 ;
        RECT  2.790 3.030 3.020 4.405 ;
        RECT  2.760 3.030 2.790 3.260 ;
        RECT  2.530 1.090 2.760 3.260 ;
        RECT  2.300 3.490 2.560 3.830 ;
        RECT  2.420 1.090 2.530 1.320 ;
        RECT  2.070 1.550 2.300 3.230 ;
        RECT  2.220 3.460 2.300 3.830 ;
        RECT  2.070 3.460 2.220 3.775 ;
        RECT  2.040 1.550 2.070 1.780 ;
        RECT  1.740 2.890 2.070 3.230 ;
        RECT  0.520 3.460 2.070 3.690 ;
        RECT  1.810 0.630 2.040 1.780 ;
        RECT  1.700 1.035 1.810 1.375 ;
        RECT  0.290 1.455 0.520 3.690 ;
        RECT  0.180 1.455 0.290 1.795 ;
        RECT  0.180 2.830 0.290 3.170 ;
    END
END BMXX1

MACRO BENCX4
    CLASS CORE ;
    FOREIGN BENCX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  27.580 1.345 27.695 1.575 ;
        RECT  27.580 2.625 27.690 2.855 ;
        RECT  27.200 1.345 27.580 2.855 ;
        RECT  23.275 1.345 27.200 1.575 ;
        RECT  23.265 2.625 27.200 2.855 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  39.975 1.820 40.120 3.220 ;
        RECT  39.970 1.820 39.975 3.240 ;
        RECT  39.740 1.515 39.970 3.240 ;
        RECT  34.950 1.515 39.740 1.745 ;
        RECT  34.940 3.010 39.740 3.240 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.790 4.005 28.985 4.235 ;
        RECT  20.560 4.005 20.790 4.410 ;
        RECT  16.925 4.180 20.560 4.410 ;
        RECT  16.695 4.005 16.925 4.410 ;
        RECT  12.325 4.005 16.695 4.235 ;
        RECT  12.095 4.005 12.325 4.315 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.510 3.430 16.740 3.775 ;
        RECT  12.805 3.545 16.510 3.775 ;
        RECT  12.575 3.075 12.805 3.775 ;
        RECT  9.455 3.105 12.575 3.335 ;
        RECT  9.245 2.940 9.455 3.335 ;
        RECT  9.015 2.560 9.245 3.335 ;
        RECT  7.405 2.965 9.015 3.195 ;
        RECT  7.175 2.580 7.405 3.195 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.400 0.635 13.560 1.955 ;
        RECT  13.330 0.635 13.400 2.385 ;
        RECT  12.640 0.635 13.330 0.865 ;
        RECT  13.170 1.725 13.330 2.385 ;
        RECT  12.410 0.635 12.640 1.035 ;
        RECT  10.970 0.805 12.410 1.035 ;
        RECT  10.740 0.805 10.970 2.050 ;
        RECT  8.365 1.820 10.740 2.050 ;
        RECT  8.135 1.820 8.365 2.635 ;
        RECT  8.060 1.955 8.135 2.635 ;
        RECT  7.550 1.955 8.060 2.185 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 1.390 5.085 1.730 ;
        RECT  1.185 2.740 5.085 3.080 ;
        RECT  1.180 1.390 1.185 3.080 ;
        RECT  0.900 1.390 1.180 3.220 ;
        RECT  0.800 1.820 0.900 3.220 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  40.050 -0.400 40.260 0.400 ;
        RECT  39.710 -0.400 40.050 1.110 ;
        RECT  38.690 -0.400 39.710 0.400 ;
        RECT  38.350 -0.400 38.690 1.110 ;
        RECT  37.330 -0.400 38.350 0.400 ;
        RECT  36.990 -0.400 37.330 1.110 ;
        RECT  35.970 -0.400 36.990 0.400 ;
        RECT  35.630 -0.400 35.970 1.110 ;
        RECT  34.610 -0.400 35.630 0.400 ;
        RECT  34.270 -0.400 34.610 1.110 ;
        RECT  33.135 -0.400 34.270 0.400 ;
        RECT  33.135 0.770 33.285 1.110 ;
        RECT  32.795 -0.400 33.135 1.110 ;
        RECT  31.335 -0.400 32.795 0.400 ;
        RECT  32.475 0.770 32.795 1.110 ;
        RECT  30.995 -0.400 31.335 0.575 ;
        RECT  28.375 -0.400 30.995 0.400 ;
        RECT  28.035 -0.400 28.375 0.575 ;
        RECT  27.015 -0.400 28.035 0.400 ;
        RECT  26.675 -0.400 27.015 0.575 ;
        RECT  25.655 -0.400 26.675 0.400 ;
        RECT  25.315 -0.400 25.655 0.575 ;
        RECT  24.295 -0.400 25.315 0.400 ;
        RECT  23.955 -0.400 24.295 0.575 ;
        RECT  22.935 -0.400 23.955 0.400 ;
        RECT  22.595 -0.400 22.935 0.575 ;
        RECT  21.575 -0.400 22.595 0.400 ;
        RECT  21.235 -0.400 21.575 0.575 ;
        RECT  15.895 -0.400 21.235 0.400 ;
        RECT  15.605 -0.400 15.895 0.575 ;
        RECT  15.605 0.980 15.895 1.320 ;
        RECT  15.375 -0.400 15.605 1.320 ;
        RECT  15.085 -0.400 15.375 0.575 ;
        RECT  15.085 0.980 15.375 1.320 ;
        RECT  12.180 -0.400 15.085 0.400 ;
        RECT  11.840 -0.400 12.180 0.575 ;
        RECT  8.840 -0.400 11.840 0.400 ;
        RECT  8.500 -0.400 8.840 0.575 ;
        RECT  7.225 -0.400 8.500 0.400 ;
        RECT  6.885 -0.400 7.225 0.950 ;
        RECT  5.725 -0.400 6.885 0.400 ;
        RECT  5.385 -0.400 5.725 0.950 ;
        RECT  4.445 -0.400 5.385 0.400 ;
        RECT  4.105 -0.400 4.445 0.950 ;
        RECT  3.165 -0.400 4.105 0.400 ;
        RECT  2.825 -0.400 3.165 0.950 ;
        RECT  1.880 -0.400 2.825 0.400 ;
        RECT  1.540 -0.400 1.880 0.950 ;
        RECT  0.600 -0.400 1.540 0.400 ;
        RECT  0.260 -0.400 0.600 0.950 ;
        RECT  0.000 -0.400 0.260 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  40.045 4.640 40.260 5.440 ;
        RECT  39.705 3.775 40.045 5.440 ;
        RECT  38.685 4.640 39.705 5.440 ;
        RECT  38.345 3.775 38.685 5.440 ;
        RECT  37.325 4.640 38.345 5.440 ;
        RECT  36.985 3.775 37.325 5.440 ;
        RECT  35.965 4.640 36.985 5.440 ;
        RECT  35.625 3.775 35.965 5.440 ;
        RECT  34.600 4.640 35.625 5.440 ;
        RECT  34.260 3.775 34.600 5.440 ;
        RECT  33.240 4.640 34.260 5.440 ;
        RECT  32.900 3.825 33.240 5.440 ;
        RECT  30.285 4.640 32.900 5.440 ;
        RECT  29.945 3.825 30.285 5.440 ;
        RECT  28.370 4.640 29.945 5.440 ;
        RECT  28.030 4.465 28.370 5.440 ;
        RECT  27.010 4.640 28.030 5.440 ;
        RECT  26.670 4.465 27.010 5.440 ;
        RECT  25.650 4.640 26.670 5.440 ;
        RECT  25.310 4.465 25.650 5.440 ;
        RECT  24.290 4.640 25.310 5.440 ;
        RECT  23.950 4.465 24.290 5.440 ;
        RECT  22.925 4.640 23.950 5.440 ;
        RECT  22.585 4.465 22.925 5.440 ;
        RECT  21.565 4.640 22.585 5.440 ;
        RECT  21.225 4.465 21.565 5.440 ;
        RECT  16.465 4.640 21.225 5.440 ;
        RECT  16.125 4.465 16.465 5.440 ;
        RECT  14.855 4.640 16.125 5.440 ;
        RECT  14.515 4.465 14.855 5.440 ;
        RECT  13.230 4.640 14.515 5.440 ;
        RECT  12.890 4.465 13.230 5.440 ;
        RECT  11.515 4.640 12.890 5.440 ;
        RECT  11.285 4.005 11.515 5.440 ;
        RECT  9.710 4.640 11.285 5.440 ;
        RECT  9.370 4.465 9.710 5.440 ;
        RECT  7.060 4.640 9.370 5.440 ;
        RECT  6.720 4.465 7.060 5.440 ;
        RECT  5.725 4.640 6.720 5.440 ;
        RECT  5.385 3.850 5.725 5.440 ;
        RECT  4.445 4.640 5.385 5.440 ;
        RECT  4.105 3.850 4.445 5.440 ;
        RECT  3.165 4.640 4.105 5.440 ;
        RECT  2.825 3.850 3.165 5.440 ;
        RECT  1.880 4.640 2.825 5.440 ;
        RECT  1.540 3.850 1.880 5.440 ;
        RECT  0.600 4.640 1.540 5.440 ;
        RECT  0.260 3.850 0.600 5.440 ;
        RECT  0.000 4.640 0.260 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  34.500 2.060 38.605 2.290 ;
        RECT  34.415 1.515 34.500 2.290 ;
        RECT  34.270 1.515 34.415 3.025 ;
        RECT  33.590 1.515 34.270 1.745 ;
        RECT  34.185 2.060 34.270 3.025 ;
        RECT  33.580 2.795 34.185 3.025 ;
        RECT  33.360 2.190 33.840 2.420 ;
        RECT  33.350 1.350 33.360 2.420 ;
        RECT  33.130 1.350 33.350 3.595 ;
        RECT  29.355 1.350 33.130 1.580 ;
        RECT  33.120 2.190 33.130 3.595 ;
        RECT  31.550 3.365 33.120 3.595 ;
        RECT  32.660 1.990 32.890 2.855 ;
        RECT  30.895 2.625 32.660 2.855 ;
        RECT  30.415 0.805 32.095 1.035 ;
        RECT  31.320 3.120 31.550 4.405 ;
        RECT  29.470 3.365 31.320 3.595 ;
        RECT  30.665 1.810 30.895 3.110 ;
        RECT  28.700 1.810 30.665 2.040 ;
        RECT  29.010 2.880 30.665 3.110 ;
        RECT  28.550 2.270 30.435 2.500 ;
        RECT  30.185 0.630 30.415 1.035 ;
        RECT  29.095 0.630 30.185 0.860 ;
        RECT  29.240 3.365 29.470 4.225 ;
        RECT  28.780 2.880 29.010 3.775 ;
        RECT  20.300 3.545 28.780 3.775 ;
        RECT  28.470 0.805 28.700 2.040 ;
        RECT  28.320 2.270 28.550 3.315 ;
        RECT  21.005 0.805 28.470 1.035 ;
        RECT  21.015 3.085 28.320 3.315 ;
        RECT  22.300 1.890 26.930 2.120 ;
        RECT  22.200 1.890 22.300 2.855 ;
        RECT  22.070 1.290 22.200 2.855 ;
        RECT  21.970 1.290 22.070 2.120 ;
        RECT  21.905 2.625 22.070 2.855 ;
        RECT  20.545 1.890 21.730 2.120 ;
        RECT  20.785 2.535 21.015 3.315 ;
        RECT  20.775 0.630 21.005 1.035 ;
        RECT  20.135 2.535 20.785 2.765 ;
        RECT  16.420 0.630 20.775 0.860 ;
        RECT  20.315 1.090 20.545 2.305 ;
        RECT  17.425 1.090 20.315 1.320 ;
        RECT  19.695 2.075 20.315 2.305 ;
        RECT  20.070 3.545 20.300 3.950 ;
        RECT  19.235 1.550 20.085 1.780 ;
        RECT  17.395 3.720 20.070 3.950 ;
        RECT  19.465 2.075 19.695 3.490 ;
        RECT  17.705 3.260 19.465 3.490 ;
        RECT  19.005 1.550 19.235 3.030 ;
        RECT  17.145 1.550 19.005 1.780 ;
        RECT  17.395 2.800 19.005 3.030 ;
        RECT  16.935 2.270 18.775 2.500 ;
        RECT  17.165 2.800 17.395 3.200 ;
        RECT  17.165 3.490 17.395 3.950 ;
        RECT  16.285 2.970 17.165 3.200 ;
        RECT  16.985 3.490 17.165 3.720 ;
        RECT  16.915 1.265 17.145 1.780 ;
        RECT  16.705 2.270 16.935 2.740 ;
        RECT  16.705 1.265 16.915 1.495 ;
        RECT  14.660 2.510 16.705 2.740 ;
        RECT  16.190 0.630 16.420 2.215 ;
        RECT  16.055 2.970 16.285 3.260 ;
        RECT  14.510 1.985 16.190 2.215 ;
        RECT  15.365 3.030 16.055 3.260 ;
        RECT  14.430 2.510 14.660 3.315 ;
        RECT  14.280 0.715 14.510 2.215 ;
        RECT  13.265 3.085 14.430 3.315 ;
        RECT  14.125 1.985 14.280 2.215 ;
        RECT  13.895 1.985 14.125 2.855 ;
        RECT  13.690 2.625 13.895 2.855 ;
        RECT  13.035 2.615 13.265 3.315 ;
        RECT  12.935 1.095 13.100 1.495 ;
        RECT  12.935 2.615 13.035 2.845 ;
        RECT  12.870 1.095 12.935 2.845 ;
        RECT  12.705 1.265 12.870 2.845 ;
        RECT  11.990 2.545 12.705 2.775 ;
        RECT  11.515 1.265 11.770 1.495 ;
        RECT  11.285 1.265 11.515 2.510 ;
        RECT  11.015 2.280 11.285 2.510 ;
        RECT  10.665 2.280 11.015 2.870 ;
        RECT  9.630 2.280 10.665 2.510 ;
        RECT  9.340 0.635 10.480 0.865 ;
        RECT  6.830 1.355 10.480 1.585 ;
        RECT  8.335 3.565 10.470 3.795 ;
        RECT  9.110 0.635 9.340 1.035 ;
        RECT  7.740 0.805 9.110 1.035 ;
        RECT  8.105 3.500 8.335 4.310 ;
        RECT  6.830 3.500 8.105 3.730 ;
        RECT  6.600 1.355 6.830 3.730 ;
        RECT  6.260 2.090 6.600 2.430 ;
        RECT  6.030 1.390 6.370 1.730 ;
        RECT  6.030 2.740 6.370 3.080 ;
        RECT  6.025 1.500 6.030 1.730 ;
        RECT  6.025 2.740 6.030 2.970 ;
        RECT  5.795 1.500 6.025 2.970 ;
        RECT  5.325 2.155 5.795 2.385 ;
        RECT  4.515 2.100 5.325 2.440 ;
        RECT  3.120 2.155 4.515 2.385 ;
        RECT  2.310 2.100 3.120 2.440 ;
    END
END BENCX4

MACRO BENCX2
    CLASS CORE ;
    FOREIGN BENCX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BENCX4 ;
    SIZE 27.060 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.945 1.265 18.855 1.495 ;
        RECT  17.945 2.625 18.285 2.855 ;
        RECT  17.715 1.265 17.945 2.855 ;
        RECT  16.985 1.265 17.715 1.495 ;
        RECT  17.605 2.380 17.715 2.855 ;
        RECT  17.020 2.625 17.605 2.855 ;
        RECT  16.640 2.380 17.020 2.855 ;
        RECT  16.425 2.625 16.640 2.855 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.110 2.965 26.185 3.195 ;
        RECT  25.960 1.315 26.110 3.195 ;
        RECT  25.955 1.315 25.960 3.720 ;
        RECT  25.880 1.260 25.955 3.720 ;
        RECT  25.720 1.260 25.880 1.545 ;
        RECT  25.620 2.965 25.880 3.720 ;
        RECT  25.380 1.205 25.720 1.545 ;
        RECT  25.525 2.965 25.620 3.220 ;
        RECT  24.635 2.965 25.525 3.195 ;
        RECT  24.280 1.260 25.380 1.545 ;
        RECT  24.520 2.965 24.635 3.220 ;
        RECT  24.290 2.965 24.520 3.740 ;
        RECT  24.180 3.400 24.290 3.740 ;
        RECT  23.940 1.205 24.280 1.545 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.545 4.055 19.655 4.285 ;
        RECT  19.315 4.005 19.545 4.285 ;
        RECT  15.135 4.005 19.315 4.235 ;
        RECT  14.905 4.005 15.135 4.410 ;
        RECT  11.140 4.180 14.905 4.410 ;
        RECT  10.910 4.005 11.140 4.410 ;
        RECT  9.685 4.005 10.910 4.235 ;
        RECT  9.455 4.005 9.685 4.315 ;
        RECT  9.220 4.005 9.455 4.235 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.720 2.770 11.775 3.000 ;
        RECT  10.490 2.770 10.720 3.775 ;
        RECT  8.325 3.545 10.490 3.775 ;
        RECT  8.095 3.545 8.325 4.360 ;
        RECT  5.800 3.545 8.095 3.775 ;
        RECT  5.800 2.305 6.080 2.535 ;
        RECT  5.570 2.305 5.800 3.775 ;
        RECT  5.495 2.965 5.570 3.195 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 0.630 10.070 0.860 ;
        RECT  8.665 0.630 8.895 1.035 ;
        RECT  7.780 0.805 8.665 1.035 ;
        RECT  7.570 0.805 7.780 1.285 ;
        RECT  7.340 0.805 7.570 2.235 ;
        RECT  6.540 2.005 7.340 2.235 ;
        RECT  6.310 1.845 6.540 2.235 ;
        RECT  5.140 1.845 6.310 2.075 ;
        RECT  4.910 1.845 5.140 2.635 ;
        RECT  4.835 2.405 4.910 2.635 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 0.835 2.690 1.645 ;
        RECT  2.350 3.090 2.690 3.955 ;
        RECT  1.250 1.415 2.350 1.645 ;
        RECT  1.535 3.090 2.350 3.320 ;
        RECT  1.250 2.940 1.535 3.320 ;
        RECT  0.910 0.835 1.250 3.955 ;
        RECT  0.875 2.405 0.910 2.635 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.385 -0.400 27.060 0.400 ;
        RECT  26.155 -0.400 26.385 0.955 ;
        RECT  25.000 -0.400 26.155 0.400 ;
        RECT  24.660 -0.400 25.000 0.965 ;
        RECT  23.520 -0.400 24.660 0.400 ;
        RECT  23.180 -0.400 23.520 0.575 ;
        RECT  22.400 -0.400 23.180 0.400 ;
        RECT  22.060 -0.400 22.400 0.575 ;
        RECT  20.875 -0.400 22.060 0.400 ;
        RECT  20.535 -0.400 20.875 0.575 ;
        RECT  18.090 -0.400 20.535 0.400 ;
        RECT  17.750 -0.400 18.090 0.575 ;
        RECT  16.565 -0.400 17.750 0.400 ;
        RECT  16.225 -0.400 16.565 0.575 ;
        RECT  11.910 -0.400 16.225 0.400 ;
        RECT  11.570 -0.400 11.910 0.575 ;
        RECT  10.530 -0.400 11.570 0.400 ;
        RECT  10.300 -0.400 10.530 1.380 ;
        RECT  8.430 -0.400 10.300 0.400 ;
        RECT  10.050 1.150 10.300 1.380 ;
        RECT  8.090 -0.400 8.430 0.575 ;
        RECT  4.970 -0.400 8.090 0.400 ;
        RECT  4.630 -0.400 4.970 0.575 ;
        RECT  3.450 -0.400 4.630 0.400 ;
        RECT  3.110 -0.400 3.450 1.090 ;
        RECT  1.970 -0.400 3.110 0.400 ;
        RECT  1.630 -0.400 1.970 1.050 ;
        RECT  0.530 -0.400 1.630 0.400 ;
        RECT  0.190 -0.400 0.530 1.490 ;
        RECT  0.000 -0.400 0.190 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.625 4.640 27.060 5.440 ;
        RECT  26.395 3.550 26.625 5.440 ;
        RECT  25.240 4.640 26.395 5.440 ;
        RECT  24.900 3.550 25.240 5.440 ;
        RECT  23.760 4.640 24.900 5.440 ;
        RECT  23.420 3.430 23.760 5.440 ;
        RECT  22.160 4.640 23.420 5.440 ;
        RECT  21.820 4.465 22.160 5.440 ;
        RECT  20.280 4.640 21.820 5.440 ;
        RECT  19.940 4.465 20.280 5.440 ;
        RECT  19.085 4.640 19.940 5.440 ;
        RECT  18.745 4.465 19.085 5.440 ;
        RECT  17.525 4.640 18.745 5.440 ;
        RECT  17.185 4.465 17.525 5.440 ;
        RECT  16.005 4.640 17.185 5.440 ;
        RECT  15.665 4.465 16.005 5.440 ;
        RECT  10.680 4.640 15.665 5.440 ;
        RECT  10.340 4.465 10.680 5.440 ;
        RECT  7.795 4.640 10.340 5.440 ;
        RECT  7.565 4.005 7.795 5.440 ;
        RECT  6.290 4.640 7.565 5.440 ;
        RECT  5.950 4.465 6.290 5.440 ;
        RECT  4.930 4.640 5.950 5.440 ;
        RECT  4.590 4.465 4.930 5.440 ;
        RECT  3.410 4.640 4.590 5.440 ;
        RECT  3.070 4.020 3.410 5.440 ;
        RECT  1.970 4.640 3.070 5.440 ;
        RECT  1.630 3.550 1.970 5.440 ;
        RECT  0.530 4.640 1.630 5.440 ;
        RECT  0.190 3.550 0.530 5.440 ;
        RECT  0.000 4.640 0.190 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  24.040 2.100 24.850 2.440 ;
        RECT  23.295 2.155 24.040 2.385 ;
        RECT  23.065 1.285 23.295 3.025 ;
        RECT  22.620 1.285 23.065 1.515 ;
        RECT  22.580 2.795 23.065 3.025 ;
        RECT  22.215 2.065 22.555 2.405 ;
        RECT  21.690 2.120 22.215 2.350 ;
        RECT  21.460 1.445 21.690 3.615 ;
        RECT  21.410 0.985 21.635 1.215 ;
        RECT  20.885 1.445 21.460 1.675 ;
        RECT  19.665 3.385 21.460 3.615 ;
        RECT  21.180 0.805 21.410 1.215 ;
        RECT  20.340 2.360 21.230 2.590 ;
        RECT  20.260 0.805 21.180 1.035 ;
        RECT  20.655 1.350 20.885 1.675 ;
        RECT  19.565 1.350 20.655 1.580 ;
        RECT  20.110 1.810 20.340 3.110 ;
        RECT  20.030 0.630 20.260 1.035 ;
        RECT  19.330 1.810 20.110 2.040 ;
        RECT  19.205 2.880 20.110 3.110 ;
        RECT  19.575 0.630 20.030 0.860 ;
        RECT  18.745 2.300 19.880 2.530 ;
        RECT  19.435 3.385 19.665 3.775 ;
        RECT  19.100 0.805 19.330 2.040 ;
        RECT  18.975 2.880 19.205 3.775 ;
        RECT  15.675 0.805 19.100 1.035 ;
        RECT  14.670 3.545 18.975 3.775 ;
        RECT  18.515 2.300 18.745 3.315 ;
        RECT  14.670 3.085 18.515 3.315 ;
        RECT  15.745 1.890 16.710 2.120 ;
        RECT  15.515 1.290 15.745 2.120 ;
        RECT  15.445 0.630 15.675 1.035 ;
        RECT  15.460 1.890 15.515 2.120 ;
        RECT  15.230 1.890 15.460 2.855 ;
        RECT  12.810 0.630 15.445 0.860 ;
        RECT  14.905 2.625 15.230 2.855 ;
        RECT  14.210 1.090 14.720 1.320 ;
        RECT  14.440 2.545 14.670 3.315 ;
        RECT  14.440 3.545 14.670 3.945 ;
        RECT  11.805 3.715 14.440 3.945 ;
        RECT  13.980 1.090 14.210 3.485 ;
        RECT  13.090 1.090 13.980 1.320 ;
        RECT  12.525 3.255 13.980 3.485 ;
        RECT  13.520 1.640 13.750 3.025 ;
        RECT  12.860 1.640 13.520 1.870 ;
        RECT  12.295 2.795 13.520 3.025 ;
        RECT  12.695 2.265 13.290 2.495 ;
        RECT  12.630 1.265 12.860 1.870 ;
        RECT  12.580 0.630 12.810 1.035 ;
        RECT  12.465 2.265 12.695 2.540 ;
        RECT  12.370 1.265 12.630 1.495 ;
        RECT  11.735 0.805 12.580 1.035 ;
        RECT  10.260 2.310 12.465 2.540 ;
        RECT  12.065 2.795 12.295 3.460 ;
        RECT  11.735 1.715 12.065 1.945 ;
        RECT  11.185 3.230 12.065 3.460 ;
        RECT  11.505 0.805 11.735 1.945 ;
        RECT  11.095 1.715 11.505 1.945 ;
        RECT  10.955 3.230 11.185 3.655 ;
        RECT  10.865 0.950 11.095 1.945 ;
        RECT  9.760 1.715 10.865 1.945 ;
        RECT  10.030 2.310 10.260 3.315 ;
        RECT  8.775 3.085 10.030 3.315 ;
        RECT  9.530 1.715 9.760 2.855 ;
        RECT  9.355 1.150 9.675 1.380 ;
        RECT  9.255 2.625 9.530 2.855 ;
        RECT  9.125 1.150 9.355 1.495 ;
        RECT  8.775 1.265 9.125 1.495 ;
        RECT  8.545 1.265 8.775 3.315 ;
        RECT  8.270 3.085 8.545 3.315 ;
        RECT  8.025 1.535 8.255 2.700 ;
        RECT  7.445 2.470 8.025 2.700 ;
        RECT  7.215 2.470 7.445 3.225 ;
        RECT  7.165 2.995 7.215 3.225 ;
        RECT  6.800 2.995 7.165 3.315 ;
        RECT  7.000 1.545 7.110 1.775 ;
        RECT  6.945 0.825 7.090 1.055 ;
        RECT  4.970 4.005 7.050 4.235 ;
        RECT  6.770 1.385 7.000 1.775 ;
        RECT  6.715 0.825 6.945 1.155 ;
        RECT  6.280 2.995 6.800 3.225 ;
        RECT  4.670 1.385 6.770 1.615 ;
        RECT  5.390 0.925 6.715 1.155 ;
        RECT  4.740 3.025 4.970 4.235 ;
        RECT  3.895 3.025 4.740 3.255 ;
        RECT  4.440 1.385 4.670 2.010 ;
        RECT  3.895 1.780 4.440 2.010 ;
        RECT  4.060 0.845 4.210 1.185 ;
        RECT  3.790 3.550 4.130 4.360 ;
        RECT  3.830 0.845 4.060 1.550 ;
        RECT  3.665 1.780 3.895 3.255 ;
        RECT  3.155 1.320 3.830 1.550 ;
        RECT  3.155 3.550 3.790 3.780 ;
        RECT  3.555 1.780 3.665 2.120 ;
        RECT  2.925 1.320 3.155 3.780 ;
        RECT  2.115 2.100 2.925 2.440 ;
    END
END BENCX2

MACRO BENCX1
    CLASS CORE ;
    FOREIGN BENCX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BENCX4 ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE smic18site ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.060 1.265 14.290 2.855 ;
        RECT  13.785 1.265 14.060 1.495 ;
        RECT  13.900 2.380 14.060 2.855 ;
        RECT  13.340 2.380 13.900 2.660 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.015 1.315 20.245 3.220 ;
        RECT  19.545 1.315 20.015 1.545 ;
        RECT  19.560 2.990 20.015 3.220 ;
        RECT  19.330 2.990 19.560 3.740 ;
        RECT  19.205 1.205 19.545 1.545 ;
        RECT  19.280 3.220 19.330 3.740 ;
        RECT  19.220 3.400 19.280 3.740 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.670 4.055 15.915 4.285 ;
        RECT  15.440 4.055 15.670 4.350 ;
        RECT  14.075 4.120 15.440 4.350 ;
        RECT  13.940 4.060 14.075 4.350 ;
        RECT  13.710 4.005 13.940 4.350 ;
        RECT  12.800 4.005 13.710 4.235 ;
        RECT  12.570 4.005 12.800 4.410 ;
        RECT  9.715 4.180 12.570 4.410 ;
        RECT  9.485 4.005 9.715 4.410 ;
        RECT  7.705 4.005 9.485 4.235 ;
        RECT  7.475 4.005 7.705 4.315 ;
        RECT  6.965 4.005 7.475 4.235 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.070 2.770 10.115 3.000 ;
        RECT  8.840 2.770 9.070 3.775 ;
        RECT  6.635 3.545 8.840 3.775 ;
        RECT  6.295 3.545 6.635 3.830 ;
        RECT  4.315 3.545 6.295 3.775 ;
        RECT  4.085 2.750 4.315 3.775 ;
        RECT  3.905 2.750 4.085 3.220 ;
        RECT  3.440 2.940 3.905 3.220 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.250 0.785 7.695 1.015 ;
        RECT  7.020 0.785 7.250 1.035 ;
        RECT  5.620 0.805 7.020 1.035 ;
        RECT  5.390 0.805 5.620 2.455 ;
        RECT  3.215 2.225 5.390 2.455 ;
        RECT  2.985 2.225 3.215 2.635 ;
        RECT  2.855 2.405 2.985 2.635 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 2.740 1.200 3.080 ;
        RECT  0.820 1.460 1.160 1.800 ;
        RECT  0.875 2.740 1.145 3.195 ;
        RECT  0.860 2.740 0.875 3.080 ;
        RECT  0.555 2.740 0.860 2.970 ;
        RECT  0.800 1.540 0.820 1.800 ;
        RECT  0.555 1.570 0.800 1.800 ;
        RECT  0.325 1.570 0.555 2.970 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.265 -0.400 20.460 0.400 ;
        RECT  19.925 -0.400 20.265 0.965 ;
        RECT  18.785 -0.400 19.925 0.400 ;
        RECT  18.445 -0.400 18.785 0.575 ;
        RECT  17.625 -0.400 18.445 0.400 ;
        RECT  17.285 -0.400 17.625 0.575 ;
        RECT  16.335 -0.400 17.285 0.400 ;
        RECT  15.995 -0.400 16.335 0.575 ;
        RECT  14.885 -0.400 15.995 0.400 ;
        RECT  14.545 -0.400 14.885 0.575 ;
        RECT  13.365 -0.400 14.545 0.400 ;
        RECT  13.025 -0.400 13.365 0.575 ;
        RECT  9.005 -0.400 13.025 0.400 ;
        RECT  8.665 -0.400 9.005 0.575 ;
        RECT  6.735 -0.400 8.665 0.400 ;
        RECT  6.395 -0.400 6.735 0.575 ;
        RECT  4.660 -0.400 6.395 0.400 ;
        RECT  4.320 -0.400 4.660 0.575 ;
        RECT  3.140 -0.400 4.320 0.400 ;
        RECT  2.800 -0.400 3.140 0.575 ;
        RECT  1.840 -0.400 2.800 0.400 ;
        RECT  1.500 -0.400 1.840 0.575 ;
        RECT  0.520 -0.400 1.500 0.400 ;
        RECT  0.180 -0.400 0.520 1.050 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.280 4.640 20.460 5.440 ;
        RECT  19.940 3.595 20.280 5.440 ;
        RECT  18.800 4.640 19.940 5.440 ;
        RECT  18.460 4.465 18.800 5.440 ;
        RECT  16.485 4.640 18.460 5.440 ;
        RECT  16.145 4.465 16.485 5.440 ;
        RECT  13.480 4.640 16.145 5.440 ;
        RECT  13.140 4.465 13.480 5.440 ;
        RECT  8.915 4.640 13.140 5.440 ;
        RECT  8.575 4.465 8.915 5.440 ;
        RECT  6.065 4.640 8.575 5.440 ;
        RECT  5.835 4.005 6.065 5.440 ;
        RECT  4.465 4.640 5.835 5.440 ;
        RECT  4.125 4.465 4.465 5.440 ;
        RECT  1.880 4.640 4.125 5.440 ;
        RECT  1.540 4.465 1.880 5.440 ;
        RECT  0.520 4.640 1.540 5.440 ;
        RECT  0.180 3.470 0.520 5.440 ;
        RECT  0.000 4.640 0.180 5.440 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.965 2.100 19.305 2.440 ;
        RECT  18.335 2.155 18.965 2.385 ;
        RECT  18.105 1.210 18.335 3.225 ;
        RECT  17.885 1.210 18.105 1.440 ;
        RECT  17.805 2.995 18.105 3.225 ;
        RECT  17.575 2.100 17.875 2.440 ;
        RECT  17.550 1.600 17.575 3.690 ;
        RECT  17.345 1.600 17.550 3.980 ;
        RECT  15.765 1.600 17.345 1.830 ;
        RECT  17.320 3.460 17.345 3.980 ;
        RECT  15.670 3.460 17.320 3.690 ;
        RECT  16.255 2.060 17.115 2.290 ;
        RECT  16.290 1.140 16.965 1.370 ;
        RECT  16.060 0.805 16.290 1.370 ;
        RECT  16.025 2.060 16.255 3.215 ;
        RECT  15.760 0.805 16.060 1.035 ;
        RECT  14.755 2.060 16.025 2.290 ;
        RECT  15.210 2.985 16.025 3.215 ;
        RECT  14.750 2.525 15.795 2.755 ;
        RECT  15.535 1.350 15.765 1.830 ;
        RECT  15.530 0.630 15.760 1.035 ;
        RECT  15.440 3.460 15.670 3.810 ;
        RECT  15.265 1.350 15.535 1.580 ;
        RECT  15.245 0.630 15.530 0.860 ;
        RECT  14.980 2.985 15.210 3.775 ;
        RECT  12.340 3.545 14.980 3.775 ;
        RECT  14.525 0.805 14.755 2.290 ;
        RECT  14.520 2.525 14.750 3.315 ;
        RECT  12.800 0.805 14.525 1.035 ;
        RECT  12.340 3.085 14.520 3.315 ;
        RECT  12.805 1.890 13.830 2.120 ;
        RECT  12.805 2.625 12.915 2.855 ;
        RECT  12.575 1.890 12.805 2.855 ;
        RECT  12.570 0.630 12.800 1.035 ;
        RECT  12.340 1.890 12.575 2.120 ;
        RECT  11.085 0.630 12.570 0.860 ;
        RECT  12.110 1.115 12.340 2.120 ;
        RECT  12.110 2.525 12.340 3.315 ;
        RECT  12.110 3.545 12.340 3.945 ;
        RECT  9.945 3.715 12.110 3.945 ;
        RECT  11.650 1.090 11.880 3.485 ;
        RECT  11.500 1.090 11.650 1.405 ;
        RECT  10.805 3.255 11.650 3.485 ;
        RECT  9.985 1.175 11.500 1.405 ;
        RECT  11.190 1.640 11.420 3.025 ;
        RECT  9.670 1.640 11.190 1.870 ;
        RECT  10.575 2.795 11.190 3.025 ;
        RECT  10.730 0.630 11.085 0.945 ;
        RECT  9.720 2.100 10.880 2.330 ;
        RECT  9.465 0.715 10.730 0.945 ;
        RECT  10.345 2.795 10.575 3.460 ;
        RECT  9.530 3.230 10.345 3.460 ;
        RECT  9.490 2.100 9.720 2.540 ;
        RECT  9.440 1.320 9.670 1.870 ;
        RECT  9.300 3.230 9.530 3.655 ;
        RECT  8.610 2.310 9.490 2.540 ;
        RECT  9.235 0.715 9.465 1.035 ;
        RECT  9.225 1.320 9.440 1.550 ;
        RECT  8.985 0.805 9.235 1.035 ;
        RECT  8.985 1.850 9.205 2.080 ;
        RECT  8.755 0.805 8.985 2.080 ;
        RECT  8.295 1.850 8.755 2.080 ;
        RECT  8.380 2.310 8.610 3.315 ;
        RECT  7.580 3.085 8.380 3.315 ;
        RECT  8.150 1.315 8.295 2.080 ;
        RECT  8.065 1.315 8.150 2.855 ;
        RECT  7.905 1.315 8.065 1.545 ;
        RECT  7.920 1.850 8.065 2.855 ;
        RECT  7.810 2.625 7.920 2.855 ;
        RECT  7.350 1.315 7.580 3.315 ;
        RECT  7.205 1.315 7.350 1.545 ;
        RECT  6.525 3.060 7.350 3.290 ;
        RECT  5.850 1.270 6.080 3.280 ;
        RECT  4.645 3.050 5.850 3.280 ;
        RECT  3.340 4.005 5.265 4.235 ;
        RECT  2.500 1.765 5.160 1.995 ;
        RECT  4.875 0.805 5.105 1.330 ;
        RECT  3.560 0.805 4.875 1.035 ;
        RECT  3.205 3.450 3.340 4.235 ;
        RECT  3.110 3.060 3.205 4.235 ;
        RECT  2.975 3.060 3.110 3.680 ;
        RECT  2.500 3.060 2.975 3.290 ;
        RECT  1.670 3.525 2.640 3.755 ;
        RECT  1.670 1.305 2.600 1.535 ;
        RECT  2.270 1.765 2.500 3.290 ;
        RECT  1.930 2.100 2.270 2.440 ;
        RECT  1.440 1.305 1.670 3.755 ;
        RECT  0.790 2.100 1.440 2.440 ;
    END
END BENCX1

END LIBRARY
